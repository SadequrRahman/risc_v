* NGSPICE file created from uProcessor.ext - technology: scmos

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

.subckt uProcessor gnd vdd adrs_bus[15] adrs_bus[14] adrs_bus[13] adrs_bus[12] adrs_bus[11]
+ adrs_bus[10] adrs_bus[9] adrs_bus[8] adrs_bus[7] adrs_bus[6] adrs_bus[5] adrs_bus[4]
+ adrs_bus[3] adrs_bus[2] adrs_bus[1] adrs_bus[0] clock data_in[15] data_in[14] data_in[13]
+ data_in[12] data_in[11] data_in[10] data_in[9] data_in[8] data_in[7] data_in[6]
+ data_in[5] data_in[4] data_in[3] data_in[2] data_in[1] data_in[0] data_out[15] data_out[14]
+ data_out[13] data_out[12] data_out[11] data_out[10] data_out[9] data_out[8] data_out[7]
+ data_out[6] data_out[5] data_out[4] data_out[3] data_out[2] data_out[1] data_out[0]
+ mem_rd mem_wr reset
X_3155_ gnd gnd _3155_/Y vdd INVX1
X_2106_ _2891_/A gnd data_out[4] vdd BUFX2
X_3086_ gnd _3164_/B _3164_/C gnd _3087_/A vdd NAND3X1
X_3988_ _4166_/A _3920_/S _3988_/C gnd _3989_/A vdd OAI21X1
X_2939_ _2339_/Y gnd _2939_/Y vdd INVX1
X_4609_ _4612_/A _4195_/A gnd _4610_/C vdd NAND2X1
XSFILL44400x26100 gnd vdd FILL
XSFILL29680x100 gnd vdd FILL
XFILL71120x28100 gnd vdd FILL
X_3842_ _4297_/Q _3846_/B gnd _3842_/Y vdd NAND2X1
X_3911_ _4408_/Q _4392_/Q _3992_/B gnd _3914_/D vdd MUX2X1
X_2655_ _2593_/Y _2623_/Y _2650_/C _2655_/D gnd _2987_/B vdd AOI22X1
X_2724_ _2693_/B _2724_/B gnd _2727_/C vdd NOR2X1
X_3773_ _3773_/A _3775_/B gnd _3773_/Y vdd NAND2X1
X_4256_ _4423_/Q _4407_/Q _4252_/S gnd _4259_/D vdd MUX2X1
X_2586_ _2782_/A gnd _2586_/Y vdd INVX1
X_4187_ _4187_/A _4198_/B gnd _4187_/Y vdd NOR2X1
X_4325_ _4232_/A _4407_/CLK _4325_/D gnd vdd DFFPOSX1
XSFILL59440x42100 gnd vdd FILL
X_3207_ gnd gnd _3208_/C vdd INVX1
X_3069_ _2343_/Y gnd _3069_/Y vdd INVX1
X_3138_ gnd _3164_/B _3164_/C gnd _3139_/A vdd NAND3X1
XBUFX2_insert100 _4455_/Q gnd _2560_/B vdd BUFX2
XBUFX2_insert122 _3642_/Q gnd _4243_/C vdd BUFX2
XBUFX2_insert111 _2953_/Y gnd _3194_/C vdd BUFX2
XBUFX2_insert133 _3421_/Q gnd _3589_/A vdd BUFX2
XBUFX2_insert166 _4263_/Y gnd _4292_/B vdd BUFX2
XBUFX2_insert199 _3409_/Y gnd _2151_/A vdd BUFX2
XBUFX2_insert188 _4426_/Q gnd _2614_/C vdd BUFX2
X_2440_ _2440_/A _2443_/B gnd _2441_/A vdd NAND2X1
XBUFX2_insert155 _4444_/Q gnd _2193_/B vdd BUFX2
XBUFX2_insert177 _3625_/Q gnd _3562_/A vdd BUFX2
XBUFX2_insert144 _3649_/Y gnd _3706_/A vdd BUFX2
X_4041_ _4041_/A _4041_/B _4036_/B gnd _4041_/Y vdd MUX2X1
X_4110_ _3932_/A _4158_/B gnd _4112_/B vdd NOR2X1
X_2371_ _2371_/A _2136_/B gnd _2371_/Y vdd XOR2X1
X_3756_ _4281_/A _3767_/B _3755_/Y gnd _3756_/Y vdd OAI21X1
X_3825_ _4283_/A _3824_/B _3825_/C gnd _3825_/Y vdd AOI21X1
X_2638_ _2779_/B _2636_/Y gnd _2642_/B vdd NOR2X1
X_2569_ _2569_/A _2659_/A gnd _2573_/C vdd XNOR2X1
X_3687_ _3517_/Y gnd _3764_/A vdd INVX4
X_2707_ _2706_/B gnd _2717_/B vdd INVX1
X_4239_ _4239_/A _4240_/B _4239_/C gnd _4239_/Y vdd OAI21X1
X_4308_ _4046_/A _4298_/CLK _4308_/D gnd vdd DFFPOSX1
XSFILL29360x36100 gnd vdd FILL
X_3610_ _3557_/B _3574_/B gnd _3610_/Y vdd NAND2X1
X_4590_ _3546_/Y gnd _4592_/B vdd INVX1
X_2423_ _4061_/A _2665_/A gnd _2427_/B vdd NAND2X1
X_3472_ data_in[6] gnd _3472_/Y vdd INVX1
X_3541_ _3556_/B gnd _3541_/Y vdd INVX1
X_4024_ _4024_/A _4020_/B gnd _4024_/Y vdd NOR2X1
X_2285_ _2272_/B _2284_/Y _2282_/Y gnd _2289_/A vdd NAND3X1
X_2354_ _2560_/B _2283_/A gnd _3355_/A vdd OR2X2
XBUFX2_insert0 _4453_/Q gnd _4061_/A vdd BUFX2
X_3739_ _4312_/Q _3740_/B gnd _3739_/Y vdd NAND2X1
XSFILL14800x16100 gnd vdd FILL
X_3808_ _4377_/Q _3809_/B gnd _3808_/Y vdd NOR2X1
XSFILL29680x4100 gnd vdd FILL
XSFILL44400x34100 gnd vdd FILL
X_2972_ _2986_/A _2986_/B gnd _2972_/Y vdd AND2X2
X_4573_ _2138_/A _4436_/CLK _4518_/Y gnd vdd DFFPOSX1
X_3524_ _3524_/A _3523_/Y gnd _3524_/Y vdd NAND2X1
X_3386_ _3400_/C _3391_/A _3388_/A gnd _3410_/B vdd OAI21X1
X_3455_ _3434_/A _4593_/A gnd _3455_/Y vdd NAND2X1
X_2406_ _2406_/A _4588_/B gnd _2406_/Y vdd XNOR2X1
XSFILL59440x50100 gnd vdd FILL
X_4007_ _4005_/Y _4040_/B _4006_/Y gnd _4007_/Y vdd AOI21X1
X_2268_ _2268_/A _2266_/Y _2268_/C gnd _2268_/Y vdd OAI21X1
X_2337_ _2560_/B _2283_/A gnd _2337_/Y vdd AND2X2
X_2199_ _2199_/A _2199_/B gnd _2199_/Y vdd NAND2X1
XSFILL59920x28100 gnd vdd FILL
X_3240_ _2323_/Y _3240_/B _3292_/C gnd _3240_/Y vdd NAND3X1
XSFILL14320x28100 gnd vdd FILL
X_3171_ _3166_/Y _3171_/B gnd _3171_/Y vdd NOR2X1
X_2122_ _2124_/A _2122_/B _2121_/Y gnd _2088_/A vdd OAI21X1
X_2955_ _2969_/B _3324_/C gnd _3204_/B vdd NAND2X1
X_4556_ _4558_/B _4625_/Y _4556_/C _4556_/D gnd _4556_/Y vdd AOI22X1
X_4625_ _4621_/A _4623_/Y _4625_/C gnd _4625_/Y vdd OAI21X1
X_2886_ _2190_/A gnd _2914_/A vdd INVX1
X_3507_ data_in[11] gnd _3507_/Y vdd INVX1
X_3369_ gnd _3343_/B gnd _3369_/Y vdd NAND2X1
X_4487_ _4486_/B gnd _4488_/C vdd INVX1
X_3438_ _3437_/Y _3508_/B _3508_/C gnd _3438_/Y vdd NAND3X1
XSFILL29360x44100 gnd vdd FILL
X_2671_ _2671_/A _2662_/Y _2671_/C gnd _2671_/Y vdd NOR3X1
X_2740_ _2671_/A gnd _2740_/Y vdd INVX1
X_4410_ _3935_/A _4394_/CLK _4269_/Y gnd vdd DFFPOSX1
X_4341_ _4341_/Q _4407_/CLK _3900_/Y gnd vdd DFFPOSX1
X_3223_ _3223_/A _3223_/B gnd _3223_/Y vdd NOR2X1
X_4272_ _4412_/Q _4269_/B gnd _4273_/C vdd NOR2X1
X_3154_ gnd gnd _3156_/A vdd INVX1
X_2105_ _2706_/B gnd data_out[3] vdd BUFX2
X_3085_ _3085_/A _3007_/B _3032_/B gnd _3085_/Y vdd NAND3X1
X_2938_ _2938_/A _2938_/B gnd _2978_/A vdd NAND2X1
X_3987_ _4367_/Q _3921_/B gnd _3989_/B vdd NOR2X1
XSFILL14800x24100 gnd vdd FILL
X_2869_ _2869_/A _2869_/B _2864_/Y gnd _2870_/A vdd NAND3X1
X_4539_ _2150_/A gnd _4540_/B vdd INVX1
X_4608_ _3490_/B gnd _4608_/Y vdd INVX1
XSFILL28880x32100 gnd vdd FILL
XFILL71120x44100 gnd vdd FILL
X_2723_ _2723_/A _2723_/B _2722_/Y gnd _2723_/Y vdd OAI21X1
X_3910_ _3909_/Y _3910_/B _3909_/C _3906_/Y gnd _3915_/B vdd OAI22X1
X_3772_ _3805_/B _3703_/Y gnd _3772_/Y vdd NAND2X1
X_3841_ _3740_/A _3846_/B _3840_/Y gnd _4296_/D vdd OAI21X1
X_2585_ _2318_/B _2584_/Y gnd _2590_/A vdd NAND2X1
X_2654_ _2573_/C _2653_/Y gnd _2655_/D vdd NAND2X1
X_4324_ _4221_/A _4298_/CLK _3764_/Y gnd vdd DFFPOSX1
X_4255_ _4254_/Y _4255_/B _4254_/C _4255_/D gnd _4260_/B vdd OAI22X1
X_4186_ _4186_/A _4186_/B _4245_/S gnd _4186_/Y vdd MUX2X1
X_3206_ gnd gnd _3208_/A vdd INVX1
X_3137_ _2202_/Y _2977_/B _3032_/B gnd _3137_/Y vdd NAND3X1
X_3068_ _3049_/Y _3068_/B _3068_/C gnd _3068_/Y vdd NAND3X1
XSFILL59920x36100 gnd vdd FILL
XSFILL44880x14100 gnd vdd FILL
XBUFX2_insert167 _4263_/Y gnd _4283_/B vdd BUFX2
XBUFX2_insert101 _4455_/Q gnd _2569_/A vdd BUFX2
XBUFX2_insert145 _3649_/Y gnd _3732_/A vdd BUFX2
XBUFX2_insert112 _2953_/Y gnd _3324_/C vdd BUFX2
XBUFX2_insert123 _3563_/Y gnd _3570_/C vdd BUFX2
XBUFX2_insert156 _4444_/Q gnd _2891_/A vdd BUFX2
XBUFX2_insert134 _3421_/Q gnd _3564_/A vdd BUFX2
XBUFX2_insert178 _3625_/Q gnd _4612_/A vdd BUFX2
XBUFX2_insert189 _4426_/Q gnd _2896_/A vdd BUFX2
X_4040_ _4038_/Y _4040_/B _4039_/Y gnd _4040_/Y vdd AOI21X1
X_2370_ _2560_/B _2283_/A gnd _3375_/A vdd AND2X2
XSFILL14320x36100 gnd vdd FILL
X_3755_ _4320_/Q _3767_/B gnd _3755_/Y vdd NAND2X1
X_3824_ _4186_/B _3824_/B gnd _3825_/C vdd NOR2X1
X_3686_ _3729_/A _3685_/B _3686_/C gnd _4403_/D vdd AOI21X1
X_2706_ _2706_/A _2706_/B _2896_/A _2706_/D gnd _2706_/Y vdd AOI22X1
X_2637_ _2636_/Y _2779_/B _2637_/C _2673_/A gnd _2637_/Y vdd AOI22X1
X_2499_ _2497_/Y gnd _2500_/A vdd INVX1
X_2568_ _2659_/A _2567_/Y gnd _2650_/C vdd NAND2X1
X_4307_ _3862_/A _4373_/CLK _3863_/Y gnd vdd DFFPOSX1
X_4238_ _4238_/A _4233_/Y _4205_/S gnd _4238_/Y vdd MUX2X1
X_4169_ _3854_/A _4088_/B gnd _4171_/B vdd NOR2X1
X_3540_ _3561_/A _3540_/B gnd _3422_/A vdd NOR2X1
X_2422_ _2420_/Y _2422_/B gnd _2431_/B vdd NAND2X1
X_2353_ _2661_/A _2571_/B gnd _2353_/Y vdd OR2X2
X_3471_ _3513_/A _3513_/B _3470_/Y gnd _3474_/C vdd OAI21X1
X_4023_ _4418_/Q _3682_/A _4074_/S gnd _4026_/D vdd MUX2X1
X_2284_ _2288_/A gnd _2284_/Y vdd INVX1
XBUFX2_insert1 _4453_/Q gnd _2331_/A vdd BUFX2
XSFILL29520x12100 gnd vdd FILL
XSFILL59440x48100 gnd vdd FILL
X_3807_ _3740_/A _3809_/B _3807_/C gnd _3807_/Y vdd AOI21X1
X_3669_ _3475_/Y gnd _3752_/A vdd INVX4
X_3738_ _3704_/A _3651_/A gnd _3738_/Y vdd NAND2X1
X_2971_ _2971_/A _2970_/Y gnd _2990_/B vdd NOR2X1
X_4572_ _2135_/A _4436_/CLK _4511_/Y gnd vdd DFFPOSX1
X_3523_ _3495_/A _3522_/Y _3520_/Y gnd _3523_/Y vdd NAND3X1
X_2336_ _2560_/B _2283_/A gnd _2336_/Y vdd NOR2X1
X_3385_ _2965_/A _2965_/B gnd _3388_/A vdd NOR2X1
X_2405_ _2377_/A _4591_/B gnd _2407_/A vdd XNOR2X1
X_3454_ _3454_/A _3453_/Y gnd _3454_/Y vdd NAND2X1
X_4006_ _2110_/A _4040_/B _4206_/C gnd _4006_/Y vdd OAI21X1
X_2267_ _2574_/A _2101_/A _2256_/Y gnd _2268_/C vdd OAI21X1
X_2198_ _2198_/A _2194_/Y gnd _2199_/B vdd NOR2X1
XSFILL44880x22100 gnd vdd FILL
XSFILL14000x100 gnd vdd FILL
X_3170_ _3168_/Y _3170_/B _3169_/Y gnd _3171_/B vdd NAND3X1
X_2121_ _2124_/A _4588_/B gnd _2121_/Y vdd NAND2X1
XSFILL14320x44100 gnd vdd FILL
XCLKBUF1_insert30 clock gnd _4297_/CLK vdd CLKBUF1
X_2954_ _3324_/C _2946_/Y gnd _3204_/D vdd NAND2X1
XSFILL29520x4100 gnd vdd FILL
X_2885_ _2885_/A _2885_/B gnd _2919_/B vdd NAND2X1
X_4624_ _4621_/A _4250_/A gnd _4625_/C vdd NAND2X1
X_4555_ _4548_/C _4560_/B _4555_/C gnd _4555_/Y vdd NAND3X1
X_4486_ _4486_/A _4486_/B _4485_/Y gnd _4486_/Y vdd OAI21X1
X_3506_ _3513_/A _3513_/B _3506_/C gnd _3509_/C vdd OAI21X1
X_2319_ _2830_/B _2318_/B gnd _2320_/B vdd AND2X2
X_3299_ _3143_/A gnd gnd _3143_/D gnd _3299_/Y vdd AOI22X1
X_3368_ _3368_/A _3367_/Y gnd _3368_/Y vdd NOR2X1
X_3437_ data_in[1] gnd _3437_/Y vdd INVX1
X_2670_ _2670_/A _2670_/B _2669_/Y gnd _2671_/C vdd NAND3X1
X_4340_ _3897_/A _4298_/CLK _3898_/Y gnd vdd DFFPOSX1
X_3222_ _3220_/Y _3222_/B _3221_/Y gnd _3223_/B vdd NAND3X1
X_4271_ _3813_/A _4287_/B _4271_/C gnd _4411_/D vdd AOI21X1
X_2104_ _2104_/A gnd data_out[2] vdd BUFX2
X_3153_ _3152_/Y _3153_/B gnd _3153_/Y vdd NOR2X1
X_3084_ _2305_/Y _3090_/B _3110_/C gnd _3084_/Y vdd NAND3X1
X_2868_ _4206_/A _2868_/B gnd _2869_/B vdd NAND2X1
X_2937_ _2861_/Y _2937_/B _2936_/Y gnd _2938_/A vdd NAND3X1
X_4607_ _4612_/A _4605_/Y _4607_/C gnd _4517_/B vdd OAI21X1
X_3986_ _4351_/Q _3820_/A _3920_/S gnd _3989_/D vdd MUX2X1
X_4538_ _4538_/A _4228_/C gnd _4576_/D vdd AND2X2
X_4469_ _4469_/A _4467_/Y _4548_/C gnd _4469_/Y vdd NAND3X1
X_2799_ _2799_/A gnd _2801_/B vdd INVX1
XSFILL43440x50100 gnd vdd FILL
XSFILL14640x2100 gnd vdd FILL
XSFILL59600x16100 gnd vdd FILL
X_2722_ _2890_/A _2699_/B _2722_/C _2913_/D gnd _2722_/Y vdd OAI22X1
X_3771_ _3771_/A _3771_/B gnd _3805_/B vdd NOR2X1
X_3840_ _3840_/A _3846_/B gnd _3840_/Y vdd NAND2X1
X_2584_ _2830_/B gnd _2584_/Y vdd INVX1
X_2653_ _2592_/Y _2635_/Y _2653_/C gnd _2653_/Y vdd OAI21X1
X_4323_ _4032_/A _4373_/CLK _4323_/D gnd vdd DFFPOSX1
X_4254_ _4327_/Q _4199_/B _4254_/C gnd _4254_/Y vdd OAI21X1
X_4185_ _4183_/Y _4240_/B _4184_/Y gnd _4432_/D vdd AOI21X1
X_3205_ _3204_/Y _3205_/B gnd _3224_/A vdd NOR2X1
X_3067_ _3067_/A _3067_/B gnd _3068_/C vdd NOR2X1
X_3136_ _2311_/Y _3090_/B _3110_/C gnd _3140_/B vdd NAND3X1
X_3969_ _3969_/A _3921_/B gnd _3969_/Y vdd NOR2X1
XBUFX2_insert102 _4455_/Q gnd _2848_/A vdd BUFX2
XBUFX2_insert146 _3649_/Y gnd _3726_/A vdd BUFX2
XBUFX2_insert124 _3563_/Y gnd _3615_/C vdd BUFX2
XBUFX2_insert168 _4441_/Q gnd _2442_/A vdd BUFX2
XBUFX2_insert157 _4444_/Q gnd _2465_/B vdd BUFX2
XBUFX2_insert135 _3917_/Y gnd _3951_/B vdd BUFX2
XBUFX2_insert179 _3625_/Q gnd _4594_/A vdd BUFX2
XBUFX2_insert113 _2953_/Y gnd _3116_/C vdd BUFX2
XSFILL29040x32100 gnd vdd FILL
X_3823_ _4281_/A _3823_/B _3822_/Y gnd _3823_/Y vdd AOI21X1
XSFILL14320x52100 gnd vdd FILL
X_2636_ _2862_/A gnd _2636_/Y vdd INVX1
X_3685_ _4212_/B _3685_/B gnd _3686_/C vdd NOR2X1
X_2705_ _2899_/A gnd _2706_/D vdd INVX1
X_3754_ _3788_/A _3754_/B _3753_/Y gnd _3754_/Y vdd OAI21X1
X_4306_ _4024_/A _4417_/CLK _4306_/D gnd vdd DFFPOSX1
X_4237_ _4237_/A _4235_/Y _4199_/C _4237_/D gnd _4238_/A vdd OAI22X1
X_2567_ _2569_/A gnd _2567_/Y vdd INVX1
X_2498_ _2500_/B _2497_/Y gnd _3176_/A vdd XNOR2X1
X_4168_ _4415_/Q _3673_/A _4166_/B gnd _4171_/D vdd MUX2X1
X_3119_ _3114_/Y _3119_/B gnd _3120_/C vdd NOR2X1
X_4099_ _3921_/A _4158_/B gnd _4101_/B vdd NOR2X1
XSFILL44400x48100 gnd vdd FILL
X_2283_ _2283_/A _2560_/B gnd _2288_/A vdd XNOR2X1
X_2421_ _2421_/A _2421_/B gnd _2422_/B vdd XNOR2X1
X_2352_ _2331_/A _2330_/B gnd _3303_/A vdd OR2X2
X_3470_ _3146_/Y gnd _3470_/Y vdd INVX1
X_4022_ _4022_/A _4020_/Y _4021_/C _4022_/D gnd _4027_/B vdd OAI22X1
XBUFX2_insert2 _4453_/Q gnd _2101_/A vdd BUFX2
X_3806_ _4376_/Q _3809_/B gnd _3807_/C vdd NOR2X1
X_3737_ _3804_/A _3737_/B _3736_/Y gnd _4375_/D vdd OAI21X1
X_2619_ _2619_/A _2618_/Y gnd _2619_/Y vdd NAND2X1
X_3668_ _3717_/A _3671_/B _3668_/C gnd _3668_/Y vdd AOI21X1
X_3599_ _2965_/B _3605_/B gnd _3600_/A vdd NAND2X1
XSFILL59600x24100 gnd vdd FILL
X_2970_ _2964_/Y _3341_/B _2970_/C gnd _2970_/Y vdd OAI21X1
X_4571_ _4501_/B _4297_/CLK _4571_/D gnd vdd DFFPOSX1
X_3522_ _3521_/Y _3508_/B _3508_/C gnd _3522_/Y vdd NAND3X1
X_3453_ _3495_/A _3452_/Y _3450_/Y gnd _3453_/Y vdd NAND3X1
X_2404_ _2402_/Y _2404_/B gnd _2416_/A vdd NAND2X1
X_2266_ _2101_/A gnd _2266_/Y vdd INVX1
X_2335_ _2333_/Y _2335_/B gnd _3344_/A vdd NOR2X1
X_3384_ _3384_/A gnd _3387_/B vdd INVX1
X_4005_ _4005_/A _4000_/Y _4027_/S gnd _4005_/Y vdd MUX2X1
X_2197_ _2394_/B _2395_/A gnd _2198_/A vdd NOR2X1
X_2120_ _4476_/C gnd _2122_/B vdd INVX1
XCLKBUF1_insert31 clock gnd _4417_/CLK vdd CLKBUF1
X_4623_ _4623_/A gnd _4623_/Y vdd INVX1
X_2884_ _2884_/A _2915_/A _2916_/A _2884_/D gnd _2885_/B vdd AOI22X1
XSFILL29520x18100 gnd vdd FILL
X_2953_ _2965_/B _2941_/Y gnd _2953_/Y vdd NOR2X1
X_4554_ _4545_/Y _4547_/B _4553_/Y gnd _4555_/C vdd OAI21X1
X_4485_ _4488_/B gnd _4485_/Y vdd INVX1
X_3505_ _3505_/A gnd _3506_/C vdd INVX1
X_3436_ _3513_/A _3513_/B _3435_/Y gnd _3436_/Y vdd OAI21X1
X_2318_ _2830_/B _2318_/B gnd _2320_/A vdd NOR2X1
X_2249_ _2235_/Y _2249_/B gnd _2251_/A vdd NAND2X1
X_3298_ gnd _3240_/B _3324_/C gnd _3298_/Y vdd NAND3X1
X_3367_ _3365_/Y _3341_/B _3367_/C gnd _3367_/Y vdd OAI21X1
X_4270_ _4124_/A _4287_/B gnd _4271_/C vdd NOR2X1
X_2103_ _2849_/A gnd data_out[15] vdd BUFX2
X_3221_ _3143_/A gnd gnd _3143_/D gnd _3221_/Y vdd AOI22X1
X_3152_ _3150_/Y _3204_/B _3152_/C _3204_/D gnd _3152_/Y vdd OAI22X1
X_3083_ gnd _3343_/B gnd _3088_/A vdd NAND2X1
XSFILL59280x6100 gnd vdd FILL
X_3985_ _3985_/A _3941_/B _3984_/Y gnd _4446_/D vdd AOI21X1
X_2867_ _4028_/A gnd _2868_/B vdd INVX1
X_4606_ _4612_/A _4184_/A gnd _4607_/C vdd NAND2X1
X_2798_ _2799_/A _2798_/B _2614_/C _2797_/Y gnd _2798_/Y vdd OAI22X1
X_2936_ _2935_/Y _2920_/B gnd _2936_/Y vdd AND2X2
X_4537_ _4537_/A _4535_/Y _4537_/C gnd _4538_/A vdd OAI21X1
X_4468_ _4565_/Q _4470_/C gnd _4469_/A vdd NAND2X1
X_3419_ _3391_/A _3632_/CLK _3419_/D gnd vdd DFFPOSX1
X_4399_ _3673_/A _4394_/CLK _4399_/D gnd vdd DFFPOSX1
XSFILL44560x10100 gnd vdd FILL
XSFILL59600x32100 gnd vdd FILL
X_3770_ _3804_/A _3760_/B _3770_/C gnd _3770_/Y vdd OAI21X1
X_2652_ _2577_/Y _2652_/B _2651_/Y gnd _2653_/C vdd AOI21X1
X_2721_ _2716_/Y _2710_/Y _2720_/Y gnd _2721_/Y vdd OAI21X1
XFILL71280x12100 gnd vdd FILL
X_4322_ _4199_/A _4359_/CLK _4322_/D gnd vdd DFFPOSX1
X_4253_ _4253_/A _4198_/B gnd _4255_/B vdd NOR2X1
X_2583_ _2583_/A _2641_/A _2582_/Y gnd _2591_/B vdd NAND3X1
X_3204_ _3204_/A _3204_/B _3204_/C _3204_/D gnd _3204_/Y vdd OAI22X1
X_4184_ _4184_/A _4240_/B _4239_/C gnd _4184_/Y vdd OAI21X1
X_3066_ _3066_/A _3063_/Y _3065_/Y gnd _3067_/B vdd NAND3X1
X_3135_ gnd _3343_/B gnd _3140_/A vdd NAND2X1
X_2919_ _2914_/Y _2919_/B _2919_/C gnd _2919_/Y vdd OAI21X1
X_3968_ _4274_/A _4146_/B _3968_/S gnd _3971_/D vdd MUX2X1
X_3899_ _4341_/Q _3904_/B gnd _3899_/Y vdd NOR2X1
XSFILL14000x32100 gnd vdd FILL
XBUFX2_insert125 _3563_/Y gnd _3579_/C vdd BUFX2
XBUFX2_insert147 _4447_/Q gnd _2881_/B vdd BUFX2
XBUFX2_insert158 _4444_/Q gnd _2428_/A vdd BUFX2
XBUFX2_insert103 _4424_/Q gnd _2619_/A vdd BUFX2
XBUFX2_insert169 _4441_/Q gnd _2932_/B vdd BUFX2
XBUFX2_insert136 _3917_/Y gnd _4152_/B vdd BUFX2
XBUFX2_insert114 _2953_/Y gnd _3246_/C vdd BUFX2
X_3822_ _3997_/B _3823_/B gnd _3822_/Y vdd NOR2X1
X_3684_ _3510_/Y gnd _3729_/A vdd INVX4
XSFILL29520x26100 gnd vdd FILL
X_2635_ _2630_/Y _2635_/B _2634_/Y gnd _2635_/Y vdd AOI21X1
X_3753_ _4166_/A _3754_/B gnd _3753_/Y vdd NAND2X1
X_2704_ _2301_/B gnd _2706_/A vdd INVX1
X_4305_ _4191_/A _4417_/CLK _4305_/D gnd vdd DFFPOSX1
X_4236_ _4341_/Q _4252_/S _4199_/C gnd _4237_/A vdd OAI21X1
X_2497_ _2496_/Y _2497_/B gnd _2497_/Y vdd AND2X2
X_2566_ _2566_/A _2566_/B gnd _3358_/A vdd NAND2X1
X_4167_ _4166_/Y _4167_/B _4155_/C _4167_/D gnd _4172_/B vdd OAI22X1
X_3049_ _3048_/Y _3049_/B gnd _3049_/Y vdd NOR2X1
X_3118_ _3116_/Y _3115_/Y _3118_/C gnd _3119_/B vdd NAND3X1
X_4098_ _4345_/Q _4377_/Q _4098_/S gnd _4101_/D vdd MUX2X1
XSFILL59120x44100 gnd vdd FILL
XSFILL14640x8100 gnd vdd FILL
X_2420_ _4050_/A _2351_/B gnd _2420_/Y vdd XNOR2X1
X_4021_ _4199_/A _4074_/S _4021_/C gnd _4022_/A vdd OAI21X1
X_2282_ _2268_/Y _2281_/Y _2272_/Y gnd _2282_/Y vdd OAI21X1
X_2351_ _2351_/A _2351_/B gnd _3277_/A vdd OR2X2
XBUFX2_insert3 _4453_/Q gnd _2925_/B vdd BUFX2
X_3736_ _3726_/A _3726_/B _4253_/A gnd _3736_/Y vdd OAI21X1
X_3805_ _3651_/A _3805_/B gnd _3805_/Y vdd AND2X2
X_2549_ _2549_/A _2548_/Y gnd _3306_/A vdd XNOR2X1
X_2618_ _2713_/A gnd _2618_/Y vdd INVX1
X_3667_ _4146_/B _3671_/B gnd _3668_/C vdd NOR2X1
X_3598_ _3601_/A data_in[14] gnd _3598_/Y vdd NAND2X1
X_4219_ _4041_/A _4041_/B _4245_/S gnd _4219_/Y vdd MUX2X1
XSFILL44880x36100 gnd vdd FILL
XSFILL59600x40100 gnd vdd FILL
X_4570_ _4495_/A _4436_/CLK _4498_/Y gnd vdd DFFPOSX1
X_2403_ _4028_/A _4206_/A gnd _2404_/B vdd XNOR2X1
X_3521_ data_in[13] gnd _3521_/Y vdd INVX1
X_3383_ _2986_/A _3382_/Y gnd _3384_/A vdd NOR2X1
X_3452_ _3451_/Y _3508_/B _3508_/C gnd _3452_/Y vdd NAND3X1
XFILL71280x20100 gnd vdd FILL
X_4004_ _4004_/A _4004_/B _4004_/C _4004_/D gnd _4005_/A vdd OAI22X1
X_2265_ _2574_/A gnd _2268_/A vdd INVX1
X_2334_ _2661_/A _2571_/B gnd _2335_/B vdd AND2X2
X_2196_ _2196_/A _2195_/B gnd _2199_/A vdd NOR2X1
X_3719_ _3752_/A _3737_/B _3719_/C gnd _3719_/Y vdd OAI21X1
X_2952_ _2952_/A gnd _2956_/C vdd INVX1
XCLKBUF1_insert32 clock gnd _4359_/CLK vdd CLKBUF1
X_4622_ _4621_/A _4620_/Y _4622_/C gnd _4549_/B vdd OAI21X1
X_4553_ _4556_/C gnd _4553_/Y vdd INVX1
X_2883_ _2418_/A gnd _2884_/D vdd INVX1
X_3366_ gnd _3340_/B gnd _3367_/C vdd NAND2X1
X_4484_ _4484_/A _4483_/Y _4557_/C gnd _4568_/D vdd AOI21X1
XSFILL14480x12100 gnd vdd FILL
X_3435_ _3435_/A gnd _3435_/Y vdd INVX1
X_3504_ _3422_/B _4614_/A gnd _3504_/Y vdd NAND2X1
X_2248_ _2245_/Y _2247_/Y gnd _3267_/A vdd NAND2X1
X_2317_ _2317_/A _2316_/Y gnd _3188_/A vdd NOR2X1
X_3297_ _3297_/A _3141_/B gnd _3300_/B vdd NAND2X1
X_2179_ _2179_/A gnd _2179_/Y vdd INVX1
X_3220_ gnd _3194_/B _3194_/C gnd _3220_/Y vdd NAND3X1
X_2102_ _2102_/A gnd data_out[14] vdd BUFX2
X_3151_ gnd gnd _3152_/C vdd INVX1
X_3082_ _3082_/A _3082_/B gnd _3094_/B vdd NOR2X1
X_2935_ _2901_/Y _2935_/B gnd _2935_/Y vdd NOR2X1
X_3984_ _2418_/A _3951_/B _3951_/C gnd _3984_/Y vdd OAI21X1
X_2866_ _2374_/B _2865_/Y gnd _2869_/A vdd NAND2X1
X_4536_ _4558_/B _4616_/Y _2147_/A _4556_/D gnd _4537_/C vdd AOI22X1
X_4605_ _4605_/A gnd _4605_/Y vdd INVX1
X_2797_ _2104_/A gnd _2797_/Y vdd INVX1
XSFILL60080x12100 gnd vdd FILL
X_3349_ _3349_/A _3141_/B gnd _3352_/B vdd NAND2X1
X_4467_ _4460_/A _4466_/Y gnd _4467_/Y vdd NAND2X1
X_3418_ _3400_/C _3632_/CLK _3416_/Y gnd vdd DFFPOSX1
X_4398_ _4157_/B _4394_/CLK _4398_/D gnd vdd DFFPOSX1
X_2582_ _2252_/A _2252_/B gnd _2582_/Y vdd XNOR2X1
X_2651_ _2647_/Y _2577_/B _2650_/Y gnd _2651_/Y vdd OAI21X1
X_2720_ _2719_/Y _2718_/Y _2717_/Y gnd _2720_/Y vdd AOI21X1
X_4252_ _4359_/Q _3836_/A _4252_/S gnd _4255_/D vdd MUX2X1
X_4321_ _4010_/A _4417_/CLK _4321_/D gnd vdd DFFPOSX1
X_4183_ _4183_/A _4178_/Y _4205_/S gnd _4183_/Y vdd MUX2X1
X_3203_ gnd gnd _3204_/C vdd INVX1
X_3065_ _3143_/A gnd gnd _3143_/D gnd _3065_/Y vdd AOI22X1
X_3134_ _3134_/A _3133_/Y gnd _3146_/B vdd NOR2X1
X_3898_ _3764_/A _3893_/B _3898_/C gnd _3898_/Y vdd AOI21X1
X_2918_ _2916_/Y _2918_/B _2918_/C gnd _2919_/C vdd AOI21X1
X_3967_ _3966_/Y _3967_/B _3988_/C _3964_/Y gnd _3972_/B vdd OAI22X1
X_2849_ _2849_/A gnd _2926_/B vdd INVX1
X_4519_ _4574_/Q gnd _4528_/A vdd INVX2
XBUFX2_insert115 _3642_/Q gnd _4254_/C vdd BUFX2
XBUFX2_insert104 _4424_/Q gnd _2292_/B vdd BUFX2
XBUFX2_insert159 _4435_/Q gnd _4217_/A vdd BUFX2
XBUFX2_insert137 _3917_/Y gnd _4217_/B vdd BUFX2
XBUFX2_insert126 _3563_/Y gnd _3582_/C vdd BUFX2
XBUFX2_insert148 _4447_/Q gnd _2482_/B vdd BUFX2
XSFILL59120x6100 gnd vdd FILL
X_3821_ _3788_/A _3809_/B _3821_/C gnd _4383_/D vdd AOI21X1
X_3752_ _3752_/A _3740_/B _3751_/Y gnd _4318_/D vdd OAI21X1
X_3683_ _3794_/A _3683_/B _3682_/Y gnd _4402_/D vdd AOI21X1
X_2565_ _2560_/Y _2565_/B gnd _2566_/B vdd NAND2X1
X_4304_ _4002_/A _4298_/CLK _4304_/D gnd vdd DFFPOSX1
X_2634_ _2600_/A _2631_/Y _2633_/Y _2600_/Y gnd _2634_/Y vdd OAI22X1
X_2703_ _2703_/A _2703_/B gnd _2703_/Y vdd NOR2X1
X_4235_ _4057_/A _4231_/B gnd _4235_/Y vdd NOR2X1
X_2496_ _2494_/Y _2218_/B gnd _2496_/Y vdd OR2X2
XSFILL29520x42100 gnd vdd FILL
X_3117_ _3143_/A gnd gnd _3143_/D gnd _3118_/C vdd AOI22X1
X_4166_ _4166_/A _4166_/B _4155_/C gnd _4166_/Y vdd OAI21X1
XSFILL14480x20100 gnd vdd FILL
X_4097_ _4097_/A _3941_/B _4096_/Y gnd _4424_/D vdd AOI21X1
X_3048_ _3046_/Y _3204_/B _3047_/Y _3204_/D gnd _3048_/Y vdd OAI22X1
XSFILL59600x38100 gnd vdd FILL
XSFILL44560x16100 gnd vdd FILL
X_4020_ _3726_/C _4020_/B gnd _4020_/Y vdd NOR2X1
X_2281_ _2280_/Y _2254_/Y _2264_/A gnd _2281_/Y vdd AOI21X1
X_2350_ _4039_/A _4217_/A gnd _3251_/A vdd OR2X2
XFILL71280x18100 gnd vdd FILL
XBUFX2_insert4 _3772_/Y gnd _3775_/B vdd BUFX2
XSFILL44240x4100 gnd vdd FILL
X_3804_ _3804_/A _3803_/B _3804_/C gnd _3804_/Y vdd OAI21X1
X_3735_ _3902_/A _3737_/B _3734_/Y gnd _3735_/Y vdd OAI21X1
X_2548_ _2547_/Y _2548_/B gnd _2548_/Y vdd NAND2X1
X_2617_ _2752_/A _2616_/Y gnd _2617_/Y vdd NAND2X1
X_3597_ _3597_/A _3595_/Y _3615_/C gnd _3597_/Y vdd AOI21X1
X_3666_ _3666_/A gnd _3717_/A vdd INVX4
X_4218_ _4216_/Y _4217_/B _4218_/C gnd _4218_/Y vdd AOI21X1
XSFILL14000x38100 gnd vdd FILL
X_2479_ _2204_/A _2201_/B gnd _2537_/A vdd XOR2X1
X_4149_ _4149_/A _4149_/B _4170_/C _4149_/D gnd _4149_/Y vdd OAI22X1
X_3520_ _3513_/A _3513_/B _3520_/C gnd _3520_/Y vdd OAI21X1
X_2402_ _4039_/A _4217_/A gnd _2402_/Y vdd XNOR2X1
X_2333_ _2661_/A _2571_/B gnd _2333_/Y vdd NOR2X1
X_3451_ data_in[3] gnd _3451_/Y vdd INVX1
X_3382_ _2986_/B gnd _3382_/Y vdd INVX1
X_4003_ _4003_/A _4052_/S _4065_/C gnd _4004_/A vdd OAI21X1
X_2264_ _2264_/A gnd _2264_/Y vdd INVX1
X_2195_ _2191_/B _2195_/B _2194_/Y gnd _2195_/Y vdd AOI21X1
X_3649_ _3649_/A _3649_/B _3649_/C gnd _3649_/Y vdd NAND3X1
X_3718_ _3703_/B _3726_/B _4366_/Q gnd _3719_/C vdd OAI21X1
XSFILL29200x14100 gnd vdd FILL
XSFILL45040x36100 gnd vdd FILL
XCLKBUF1_insert22 clock gnd _4345_/CLK vdd CLKBUF1
X_2951_ _2433_/Y gnd _2951_/Y vdd INVX1
XCLKBUF1_insert33 clock gnd _4373_/CLK vdd CLKBUF1
X_4621_ _4621_/A _4239_/A gnd _4622_/C vdd NAND2X1
X_4552_ _4578_/Q _4556_/C _4548_/B gnd _4560_/B vdd NAND3X1
X_3503_ _3503_/A _3502_/Y gnd _3503_/Y vdd NAND2X1
X_4483_ _4558_/B _4592_/Y _4488_/A _4556_/D gnd _4483_/Y vdd AOI22X1
X_2882_ _2881_/B gnd _2884_/A vdd INVX1
X_2316_ _2218_/B _2421_/B gnd _2316_/Y vdd AND2X2
X_3296_ _3291_/Y _3296_/B _3295_/Y gnd _3301_/A vdd NAND3X1
X_3365_ gnd gnd _3365_/Y vdd INVX1
X_3434_ _3434_/A _4584_/A gnd _3434_/Y vdd NAND2X1
XSFILL29520x50100 gnd vdd FILL
X_2247_ _2249_/B _2247_/B gnd _2247_/Y vdd NAND2X1
X_2178_ _2172_/B _2168_/Y _2178_/C gnd _2278_/A vdd NAND3X1
XSFILL44560x24100 gnd vdd FILL
X_3150_ _2483_/Y gnd _3150_/Y vdd INVX1
X_2101_ _2101_/A gnd data_out[13] vdd BUFX2
XFILL71280x26100 gnd vdd FILL
X_3081_ _3081_/A _3341_/B _3081_/C gnd _3082_/B vdd OAI21X1
XSFILL44400x100 gnd vdd FILL
X_2865_ _2374_/A gnd _2865_/Y vdd INVX1
X_2934_ _2934_/A _2933_/Y gnd _2935_/B vdd NAND2X1
X_3983_ _3982_/Y _3983_/B _4027_/S gnd _3985_/A vdd MUX2X1
X_4535_ _2147_/A _4534_/Y _4548_/C gnd _4535_/Y vdd OAI21X1
X_4466_ _4470_/C gnd _4466_/Y vdd INVX1
X_2796_ _2456_/A gnd _2798_/B vdd INVX1
X_4604_ _4594_/A _4602_/Y _4603_/Y gnd _4604_/Y vdd OAI21X1
X_3348_ _3348_/A _3348_/B _3347_/Y gnd _3353_/A vdd NAND3X1
X_3279_ _3279_/A _2950_/B _3278_/Y _3201_/D gnd _3283_/B vdd OAI22X1
X_3417_ _3406_/B _3632_/CLK _3417_/D gnd vdd DFFPOSX1
X_4397_ _4146_/B _4383_/CLK _3668_/Y gnd vdd DFFPOSX1
XSFILL14000x46100 gnd vdd FILL
X_2581_ _2778_/A _2580_/Y gnd _2641_/A vdd NAND2X1
X_4320_ _4320_/Q _4407_/CLK _3756_/Y gnd vdd DFFPOSX1
X_2650_ _2650_/A _2650_/B _2650_/C gnd _2650_/Y vdd OAI21X1
X_4251_ _4251_/A _4040_/B _4250_/Y gnd _4438_/D vdd AOI21X1
X_4182_ _4181_/Y _4182_/B _4247_/C _4182_/D gnd _4183_/A vdd OAI22X1
X_3202_ _3202_/A gnd _3204_/A vdd INVX1
X_3133_ _3133_/A _3341_/B _3132_/Y gnd _3133_/Y vdd OAI21X1
XSFILL14480x18100 gnd vdd FILL
X_3064_ gnd _3240_/B _3246_/C gnd _3066_/A vdd NAND3X1
X_2848_ _2848_/A _2848_/B gnd _2848_/Y vdd NAND2X1
X_3897_ _3897_/A _3893_/B gnd _3898_/C vdd NOR2X1
X_2917_ _2915_/A _2884_/A gnd _2918_/B vdd NAND2X1
X_3966_ _3966_/A _3968_/S _3988_/C gnd _3966_/Y vdd OAI21X1
X_2779_ _2779_/A _2779_/B _2778_/Y gnd _2828_/A vdd OAI21X1
X_4449_ _4449_/Q _4451_/CLK _4449_/D gnd vdd DFFPOSX1
X_4518_ _4516_/Y _4518_/B _4557_/C gnd _4518_/Y vdd AOI21X1
XSFILL29200x22100 gnd vdd FILL
XBUFX2_insert116 _3642_/Q gnd _4155_/C vdd BUFX2
XBUFX2_insert149 _4447_/Q gnd _2312_/A vdd BUFX2
XBUFX2_insert105 _4424_/Q gnd _2429_/B vdd BUFX2
XBUFX2_insert138 _3917_/Y gnd _4130_/B vdd BUFX2
XBUFX2_insert127 _3410_/Y gnd _3518_/A vdd BUFX2
X_3682_ _3682_/A _3683_/B gnd _3682_/Y vdd NOR2X1
X_2702_ _2699_/Y _2701_/Y _2702_/C gnd _2703_/B vdd NAND3X1
X_3820_ _3820_/A _3809_/B gnd _3821_/C vdd NOR2X1
X_3751_ _3751_/A _3740_/B gnd _3751_/Y vdd NAND2X1
X_2495_ _2218_/B _2494_/Y gnd _2497_/B vdd NAND2X1
X_2564_ _2563_/Y _2554_/A _2556_/Y gnd _2565_/B vdd OAI21X1
X_2633_ _2633_/A _2633_/B _2632_/Y gnd _2633_/Y vdd OAI21X1
X_4303_ _3854_/A _4300_/CLK _4303_/D gnd vdd DFFPOSX1
X_4234_ _4056_/A _3691_/A _4252_/S gnd _4237_/D vdd MUX2X1
X_4165_ _4367_/Q _4088_/B gnd _4167_/B vdd NOR2X1
X_4096_ _2429_/B _3941_/B _4162_/C gnd _4096_/Y vdd OAI21X1
X_3116_ gnd _3194_/B _3116_/C gnd _3116_/Y vdd NAND3X1
X_3047_ gnd gnd _3047_/Y vdd INVX1
X_3949_ _3949_/A _3949_/B _3934_/C _3946_/Y gnd _3950_/A vdd OAI22X1
XSFILL44560x32100 gnd vdd FILL
X_2280_ _2280_/A _2278_/Y _2280_/C gnd _2280_/Y vdd OAI21X1
X_3803_ _4359_/Q _3803_/B gnd _3804_/C vdd NAND2X1
XBUFX2_insert5 _3772_/Y gnd _3803_/B vdd BUFX2
XFILL71280x34100 gnd vdd FILL
X_3734_ _3732_/A _3726_/B _4064_/A gnd _3734_/Y vdd OAI21X1
X_3665_ _4273_/A _3671_/B _3664_/Y gnd _3665_/Y vdd AOI21X1
X_2616_ _2711_/A gnd _2616_/Y vdd INVX1
X_4217_ _4217_/A _4217_/B _4239_/C gnd _4218_/C vdd OAI21X1
X_2547_ _2330_/B _2544_/Y gnd _2547_/Y vdd NAND2X1
X_3596_ _2986_/A _3605_/B gnd _3597_/A vdd NAND2X1
X_2478_ _2201_/B _2478_/B gnd _2491_/B vdd NOR2X1
X_4079_ _3870_/A _4002_/B gnd _4079_/Y vdd NOR2X1
X_4148_ _3970_/A _4153_/S _4155_/C gnd _4149_/A vdd OAI21X1
X_2332_ _2330_/Y _2332_/B gnd _3318_/A vdd NOR2X1
X_2401_ _2385_/Y _2401_/B gnd _2984_/A vdd NOR2X1
X_3381_ _3601_/A gnd _3416_/A vdd INVX1
X_3450_ _3513_/A _3513_/B _3449_/Y gnd _3450_/Y vdd OAI21X1
X_4002_ _4002_/A _4002_/B gnd _4004_/B vdd NOR2X1
X_2263_ _2259_/B _2263_/B gnd _2264_/A vdd NAND2X1
X_2194_ _2394_/B _2395_/A gnd _2194_/Y vdd AND2X2
XSFILL29520x48100 gnd vdd FILL
XSFILL14480x26100 gnd vdd FILL
X_3579_ _3579_/A _3579_/B _3579_/C gnd _3579_/Y vdd AOI21X1
X_3717_ _3717_/A _3737_/B _3716_/Y gnd _4365_/D vdd OAI21X1
X_3648_ _3699_/A _3771_/A gnd _3651_/B vdd NOR2X1
XSFILL44080x44100 gnd vdd FILL
XCLKBUF1_insert23 clock gnd _4436_/CLK vdd CLKBUF1
X_4620_ _4620_/A gnd _4620_/Y vdd INVX1
X_2881_ _2879_/Y _2881_/B _2881_/C _2881_/D gnd _2885_/A vdd AOI22X1
XCLKBUF1_insert34 clock gnd _4383_/CLK vdd CLKBUF1
XSFILL14160x100 gnd vdd FILL
X_2950_ _2939_/Y _2950_/B _2950_/C _3201_/D gnd _2950_/Y vdd OAI22X1
X_4551_ _4551_/A _4228_/C gnd _4551_/Y vdd AND2X2
X_4482_ _4548_/C _4482_/B _4493_/B gnd _4484_/A vdd NAND3X1
X_3433_ _3422_/Y _3433_/B gnd _3433_/Y vdd NAND2X1
X_3502_ _3495_/A _3501_/Y _3499_/Y gnd _3502_/Y vdd NAND3X1
X_2246_ _2233_/Y _2236_/Y gnd _2247_/B vdd NOR2X1
X_2315_ _2421_/A _2421_/B gnd _2317_/A vdd NOR2X1
X_3295_ _3294_/Y _3295_/B gnd _3295_/Y vdd AND2X2
X_3364_ _3362_/Y _3130_/B _3364_/C _3130_/D gnd _3368_/A vdd OAI22X1
X_2177_ _2177_/A _2178_/C gnd _2177_/Y vdd XNOR2X1
XSFILL60080x26100 gnd vdd FILL
XSFILL14960x22100 gnd vdd FILL
XSFILL44560x40100 gnd vdd FILL
X_2100_ _2100_/A gnd data_out[12] vdd BUFX2
X_3080_ gnd _3340_/B gnd _3081_/C vdd NAND2X1
X_3982_ _3982_/A _3980_/Y _3982_/C _3982_/D gnd _3982_/Y vdd OAI22X1
X_2864_ _2921_/B _2829_/B _2863_/Y _2673_/A gnd _2864_/Y vdd AOI22X1
XFILL71280x42100 gnd vdd FILL
X_2933_ _2713_/A _2292_/B gnd _2933_/Y vdd XNOR2X1
X_2795_ _2841_/A _2794_/Y _2795_/C gnd _2795_/Y vdd OAI21X1
X_4603_ _4586_/A _2136_/B gnd _4603_/Y vdd NAND2X1
X_4534_ _4528_/A _4534_/B _4528_/B gnd _4534_/Y vdd NOR3X1
X_4465_ _4465_/A _4460_/Y _4557_/C gnd _4465_/Y vdd AOI21X1
X_3416_ _3416_/A _3417_/D gnd _3416_/Y vdd NOR2X1
X_4396_ _4135_/B _4300_/CLK _3665_/Y gnd vdd DFFPOSX1
X_2229_ _2222_/Y _2223_/Y _2229_/C gnd _2229_/Y vdd OAI21X1
X_3347_ _3346_/Y _3347_/B gnd _3347_/Y vdd AND2X2
X_3278_ gnd gnd _3278_/Y vdd INVX1
X_2580_ _2098_/A gnd _2580_/Y vdd INVX1
X_4250_ _4250_/A _4217_/B _4239_/C gnd _4250_/Y vdd OAI21X1
X_4181_ _4003_/A _4245_/S _4247_/C gnd _4181_/Y vdd OAI21X1
X_3201_ _3201_/A _2950_/B _3201_/C _3201_/D gnd _3205_/B vdd OAI22X1
X_3063_ _2358_/Y _3141_/B gnd _3063_/Y vdd NAND2X1
X_3132_ gnd _3340_/B gnd _3132_/Y vdd NAND2X1
X_3965_ _4365_/Q _3921_/B gnd _3967_/B vdd NOR2X1
X_2778_ _2778_/A _2776_/D gnd _2778_/Y vdd NAND2X1
X_2847_ _2762_/A gnd _2848_/B vdd INVX1
X_3896_ _3729_/A _3896_/B _3895_/Y gnd _3896_/Y vdd AOI21X1
XSFILL14480x34100 gnd vdd FILL
X_2916_ _2916_/A _2884_/D gnd _2916_/Y vdd NOR2X1
X_4448_ _4448_/Q _4451_/CLK _4007_/Y gnd vdd DFFPOSX1
X_4379_ _4379_/Q _4373_/CLK _3813_/Y gnd vdd DFFPOSX1
X_4517_ _4558_/B _4517_/B _2138_/A _4556_/D gnd _4518_/B vdd AOI22X1
XBUFX2_insert117 _3642_/Q gnd _4111_/C vdd BUFX2
XBUFX2_insert106 _4424_/Q gnd _2433_/A vdd BUFX2
XBUFX2_insert139 _3917_/Y gnd _3941_/B vdd BUFX2
XBUFX2_insert128 _3410_/Y gnd _3532_/A vdd BUFX2
X_3681_ _3503_/Y gnd _3794_/A vdd INVX4
X_3750_ _3717_/A _3754_/B _3749_/Y gnd _3750_/Y vdd OAI21X1
X_2632_ _2890_/A _2604_/Y _2606_/C _2913_/D gnd _2632_/Y vdd OAI22X1
X_2701_ _2913_/D _2722_/C gnd _2701_/Y vdd NAND2X1
XSFILL44240x12100 gnd vdd FILL
X_4233_ _4233_/A _4231_/Y _4199_/C _4233_/D gnd _4233_/Y vdd OAI22X1
X_2494_ _2782_/A gnd _2494_/Y vdd INVX1
X_2563_ _2553_/Y gnd _2563_/Y vdd INVX1
X_4302_ _4158_/A _4394_/CLK _4302_/D gnd vdd DFFPOSX1
X_4164_ _4351_/Q _3820_/A _4153_/S gnd _4167_/D vdd MUX2X1
X_3046_ _2453_/Y gnd _3046_/Y vdd INVX1
X_4095_ _4095_/A _4095_/B _4205_/S gnd _4097_/A vdd MUX2X1
X_3115_ _2360_/Y _3141_/B gnd _3115_/Y vdd NAND2X1
X_3948_ _3948_/A _4036_/B _3934_/C gnd _3949_/A vdd OAI21X1
XSFILL29680x10100 gnd vdd FILL
X_3879_ _3948_/A _3879_/B gnd _3879_/Y vdd NOR2X1
XBUFX2_insert6 _3772_/Y gnd _3786_/B vdd BUFX2
X_3802_ _3902_/A _3802_/B _3802_/C gnd _3802_/Y vdd OAI21X1
XFILL71280x50100 gnd vdd FILL
X_3733_ _3692_/A _3737_/B _3732_/Y gnd _3733_/Y vdd OAI21X1
X_2615_ _2615_/A _2614_/Y gnd _2622_/C vdd NAND2X1
X_3664_ _4135_/B _3671_/B gnd _3664_/Y vdd NOR2X1
X_3595_ _3601_/A data_in[13] gnd _3595_/Y vdd NAND2X1
X_4216_ _4215_/Y _4211_/Y _4205_/S gnd _4216_/Y vdd MUX2X1
X_2546_ _2545_/Y gnd _2548_/B vdd INVX1
X_2477_ _2204_/A gnd _2478_/B vdd INVX1
X_4147_ _3969_/A _4088_/B gnd _4149_/B vdd NOR2X1
X_4078_ _4423_/Q _4407_/Q _4074_/S gnd _4081_/D vdd MUX2X1
X_3029_ _3027_/Y _3341_/B _3029_/C gnd _3029_/Y vdd OAI21X1
X_2400_ _2400_/A _2391_/Y _2400_/C gnd _2401_/B vdd NAND3X1
XBUFX2_insert90 _3644_/Q gnd _3992_/B vdd BUFX2
X_4001_ _4416_/Q _4400_/Q _4012_/S gnd _4004_/D vdd MUX2X1
X_2331_ _2331_/A _2574_/A gnd _2332_/B vdd AND2X2
X_2262_ _2262_/A _2263_/B gnd _3319_/A vdd XNOR2X1
X_3380_ _3380_/A _3368_/Y _3380_/C gnd _3533_/A vdd NAND3X1
X_2193_ _2892_/A _2193_/B gnd _2195_/B vdd AND2X2
X_3716_ _3706_/A _3726_/B _4365_/Q gnd _3716_/Y vdd OAI21X1
XSFILL14480x42100 gnd vdd FILL
X_2529_ _2529_/A _2500_/B _2528_/Y gnd _2529_/Y vdd OAI21X1
X_3578_ _3564_/A data_in[6] gnd _3579_/B vdd NAND2X1
X_3647_ _3433_/Y gnd _3740_/A vdd INVX4
XSFILL59920x2100 gnd vdd FILL
XSFILL13680x100 gnd vdd FILL
XCLKBUF1_insert35 clock gnd _4451_/CLK vdd CLKBUF1
X_2880_ _2880_/A gnd _2881_/C vdd INVX1
XCLKBUF1_insert24 clock gnd _3632_/CLK vdd CLKBUF1
X_4550_ _4548_/Y _4547_/Y _4549_/Y gnd _4551_/A vdd OAI21X1
X_3363_ gnd gnd _3364_/C vdd INVX1
X_4481_ _4481_/A gnd _4493_/B vdd INVX1
X_3501_ _3500_/Y _3508_/B _3508_/C gnd _3501_/Y vdd NAND3X1
X_3432_ _3495_/A _3431_/Y _3427_/Y gnd _3433_/B vdd NAND3X1
XSFILL44240x20100 gnd vdd FILL
X_2245_ _2233_/Y _2236_/Y _2244_/Y gnd _2245_/Y vdd OAI21X1
X_3294_ gnd _3294_/B _3268_/C gnd _3294_/Y vdd NAND3X1
X_2176_ _2179_/A _2180_/C gnd _2178_/C vdd NOR2X1
X_2314_ _2314_/A _2313_/Y gnd _2314_/Y vdd NOR2X1
XSFILL59760x14100 gnd vdd FILL
XSFILL29840x6100 gnd vdd FILL
X_2932_ _2392_/B _2932_/B gnd _2934_/A vdd XNOR2X1
X_3981_ _4334_/Q _3992_/B _3909_/C gnd _3982_/A vdd OAI21X1
X_2863_ _2676_/A gnd _2863_/Y vdd INVX1
X_4533_ _4540_/A _4540_/C gnd _4537_/A vdd NOR2X1
X_2794_ _2794_/A _2794_/B gnd _2794_/Y vdd NOR2X1
X_4602_ _4602_/A gnd _4602_/Y vdd INVX1
X_3346_ gnd _3346_/B _3346_/C gnd _3346_/Y vdd NAND3X1
X_4395_ _4124_/B _4436_/CLK _4395_/D gnd vdd DFFPOSX1
X_4464_ _4558_/B _4583_/Y _4565_/Q _4556_/D gnd _4465_/A vdd AOI22X1
X_3415_ _3415_/A gnd _3420_/D vdd INVX1
X_2228_ _2228_/A _2786_/A _2219_/B gnd _2229_/C vdd OAI21X1
X_2159_ _2159_/A gnd _2159_/Y vdd INVX1
X_3277_ _3277_/A gnd _3279_/A vdd INVX1
XSFILL15120x22100 gnd vdd FILL
X_4180_ _4002_/A _4180_/B gnd _4182_/B vdd NOR2X1
X_3200_ gnd gnd _3201_/C vdd INVX1
X_3062_ _3057_/Y _3062_/B _3061_/Y gnd _3067_/A vdd NAND3X1
X_3131_ gnd gnd _3133_/A vdd INVX1
X_3895_ _4214_/A _3904_/B gnd _3895_/Y vdd NOR2X1
X_2915_ _2915_/A _2884_/A gnd _2918_/C vdd NOR2X1
X_3964_ _4142_/A _3816_/A _3968_/S gnd _3964_/Y vdd MUX2X1
X_2777_ _2862_/A gnd _2779_/A vdd INVX1
XSFILL14480x50100 gnd vdd FILL
X_2846_ _2761_/A _2846_/B gnd _2846_/Y vdd NAND2X1
X_4516_ _4548_/C _4516_/B _4528_/B gnd _4516_/Y vdd NAND3X1
X_3329_ _2353_/Y gnd _3331_/A vdd INVX1
X_4378_ _4378_/Q _4373_/CLK _3811_/Y gnd vdd DFFPOSX1
X_4447_ _4447_/Q _4431_/CLK _4447_/D gnd vdd DFFPOSX1
XBUFX2_insert107 _4452_/Q gnd _2100_/A vdd BUFX2
XBUFX2_insert129 _3410_/Y gnd _3422_/B vdd BUFX2
XBUFX2_insert118 _3642_/Q gnd _4101_/C vdd BUFX2
XFILL71280x6100 gnd vdd FILL
XSFILL14640x10100 gnd vdd FILL
X_3680_ _4283_/A _3680_/B _3679_/Y gnd _4401_/D vdd AOI21X1
X_2562_ _2556_/Y _2562_/B _2559_/Y gnd _2566_/A vdd NAND3X1
X_2631_ _2482_/B _2594_/Y gnd _2631_/Y vdd NOR2X1
X_2700_ _2891_/A gnd _2722_/C vdd INVX1
XFILL71280x48100 gnd vdd FILL
X_4232_ _4232_/A _4252_/S _4199_/C gnd _4233_/A vdd OAI21X1
X_2493_ _2474_/D _2493_/B _2541_/A gnd _2500_/B vdd AOI21X1
X_4301_ _3969_/A _4300_/CLK _3851_/Y gnd vdd DFFPOSX1
X_4163_ _4163_/A _4130_/B _4162_/Y gnd _4430_/D vdd AOI21X1
X_3045_ _3043_/Y _2950_/B _3045_/C _3201_/D gnd _3049_/B vdd OAI22X1
X_4094_ _4094_/A _4092_/Y _4101_/C _4094_/D gnd _4095_/A vdd OAI22X1
X_3114_ _3114_/A _3110_/Y _3113_/Y gnd _3114_/Y vdd NAND3X1
X_3878_ _3811_/A _3896_/B _3878_/C gnd _4330_/D vdd AOI21X1
X_3947_ _3947_/A _3932_/B gnd _3949_/B vdd NOR2X1
X_2829_ _2779_/A _2829_/B _2776_/Y gnd _2831_/C vdd OAI21X1
XBUFX2_insert7 _3772_/Y gnd _3792_/B vdd BUFX2
X_3732_ _3732_/A _3726_/B _4231_/A gnd _3732_/Y vdd OAI21X1
X_3801_ _4241_/A _3803_/B gnd _3802_/C vdd NAND2X1
X_2545_ _2330_/B _2544_/Y gnd _2545_/Y vdd NOR2X1
X_2614_ _2612_/Y _2799_/A _2614_/C _2613_/Y gnd _2614_/Y vdd AOI22X1
X_3594_ _3593_/Y _3594_/B _3570_/C gnd _3634_/D vdd AOI21X1
X_3663_ _3461_/Y gnd _4273_/A vdd INVX4
X_4215_ _4215_/A _4215_/B _4243_/C _4212_/Y gnd _4215_/Y vdd OAI22X1
X_2476_ _2476_/A _2475_/Y gnd _2476_/Y vdd XNOR2X1
X_4146_ _4274_/A _4146_/B _4153_/S gnd _4149_/D vdd MUX2X1
X_4077_ _4077_/A _4075_/Y _4021_/C _4077_/D gnd _4077_/Y vdd OAI22X1
X_3028_ gnd _3340_/B gnd _3029_/C vdd NAND2X1
XSFILL29200x44100 gnd vdd FILL
XBUFX2_insert80 _4433_/Q gnd _2228_/A vdd BUFX2
XBUFX2_insert91 _3644_/Q gnd _4074_/S vdd BUFX2
X_4000_ _4000_/A _3998_/Y _4065_/C _3997_/Y gnd _4000_/Y vdd OAI22X1
X_2330_ _2331_/A _2330_/B gnd _2330_/Y vdd NOR2X1
X_2261_ _2330_/B _2331_/A gnd _2263_/B vdd XOR2X1
X_2192_ _2192_/A _2191_/Y gnd _2192_/Y vdd XNOR2X1
XBUFX2_insert290 _4428_/Q gnd _2187_/A vdd BUFX2
X_3715_ _4273_/A _3737_/B _3715_/C gnd _4364_/D vdd OAI21X1
X_2528_ _2528_/A _2507_/Y _2528_/C gnd _2528_/Y vdd AOI21X1
X_3646_ _3905_/A _4300_/CLK _3646_/D gnd vdd DFFPOSX1
X_3577_ _4170_/C _3574_/B gnd _3579_/A vdd NAND2X1
XSFILL29680x16100 gnd vdd FILL
X_2459_ _2445_/A _2459_/B _2539_/B gnd _2474_/D vdd OAI21X1
X_4129_ _4591_/B _4130_/B _4228_/C gnd _4129_/Y vdd OAI21X1
XSFILL28720x32100 gnd vdd FILL
XSFILL59280x34100 gnd vdd FILL
XCLKBUF1_insert25 clock gnd _4298_/CLK vdd CLKBUF1
X_3500_ data_in[10] gnd _3500_/Y vdd INVX1
X_3362_ gnd gnd _3362_/Y vdd INVX1
X_4480_ _4486_/A _4486_/B gnd _4481_/A vdd NOR2X1
X_3431_ _3428_/Y _3508_/B _3508_/C gnd _3431_/Y vdd NAND3X1
X_2313_ _2312_/A _2346_/B gnd _2313_/Y vdd AND2X2
X_2244_ _2249_/B gnd _2244_/Y vdd INVX1
X_3293_ _3293_/A _3345_/B _3267_/C gnd _3295_/B vdd NAND3X1
X_2175_ _2609_/A _2706_/B gnd _2179_/A vdd NOR2X1
XSFILL44720x14100 gnd vdd FILL
X_3629_ _3545_/A _3632_/CLK _3629_/D gnd vdd DFFPOSX1
XSFILL59760x30100 gnd vdd FILL
X_2931_ _2878_/A _2877_/Y gnd _2937_/B vdd AND2X2
X_3980_ _4158_/A _3943_/B gnd _3980_/Y vdd NOR2X1
X_2862_ _2862_/A gnd _2921_/B vdd INVX1
X_4532_ _2147_/A gnd _4540_/A vdd INVX1
X_4463_ _4458_/Y _4462_/B gnd _4556_/D vdd NOR2X1
X_2793_ _2619_/A gnd _2794_/B vdd INVX1
X_4601_ _4586_/A _4601_/B _4600_/Y gnd _4601_/Y vdd OAI21X1
X_3345_ _3345_/A _3345_/B _3188_/B gnd _3347_/B vdd NAND3X1
X_3276_ _3276_/A _3276_/B _3275_/Y gnd _3505_/A vdd NAND3X1
X_4394_ _3935_/B _4394_/CLK _3659_/Y gnd vdd DFFPOSX1
X_3414_ _3391_/A _3406_/B _3649_/A gnd _3415_/A vdd OAI21X1
XSFILL14480x48100 gnd vdd FILL
X_2227_ _2227_/A _2227_/B gnd _3215_/A vdd XOR2X1
X_2158_ _2158_/A _2158_/B _2157_/Y gnd _2158_/Y vdd OAI21X1
X_2089_ _2089_/A gnd adrs_bus[3] vdd BUFX2
XSFILL29200x52100 gnd vdd FILL
X_3130_ _3130_/A _3130_/B _3129_/Y _3130_/D gnd _3134_/A vdd OAI22X1
XSFILL44240x26100 gnd vdd FILL
X_3061_ _3061_/A _3059_/Y gnd _3061_/Y vdd AND2X2
X_3894_ _3794_/A _3904_/B _3893_/Y gnd _4338_/D vdd AOI21X1
X_2845_ _2762_/C gnd _2846_/B vdd INVX1
X_2914_ _2914_/A _2190_/B _2913_/Y gnd _2914_/Y vdd OAI21X1
X_3963_ _3963_/A _4152_/B _3962_/Y gnd _4444_/D vdd AOI21X1
X_2776_ _2862_/A _2776_/B _2676_/A _2776_/D gnd _2776_/Y vdd OAI22X1
X_4515_ _2135_/A _2138_/A _4514_/Y gnd _4528_/B vdd NAND3X1
X_4446_ _4446_/Q _4431_/CLK _4446_/D gnd vdd DFFPOSX1
X_3259_ gnd gnd _3260_/C vdd INVX1
X_3328_ _3328_/A _3316_/Y _3328_/C gnd _3519_/A vdd NAND3X1
XSFILL29680x24100 gnd vdd FILL
X_4377_ _4377_/Q _4345_/CLK _3809_/Y gnd vdd DFFPOSX1
XBUFX2_insert108 _4452_/Q gnd _2351_/A vdd BUFX2
XBUFX2_insert119 _3642_/Q gnd _4170_/C vdd BUFX2
XSFILL59280x42100 gnd vdd FILL
XSFILL29360x6100 gnd vdd FILL
X_2561_ _2560_/Y gnd _2562_/B vdd INVX1
X_2630_ _2625_/Y _2622_/C _2629_/Y gnd _2630_/Y vdd OAI21X1
X_2492_ _2486_/Y _2492_/B _2492_/C gnd _2541_/A vdd OAI21X1
X_4300_ _4300_/Q _4300_/CLK _3849_/Y gnd vdd DFFPOSX1
X_4231_ _4231_/A _4231_/B gnd _4231_/Y vdd NOR2X1
X_4162_ _4600_/B _4130_/B _4162_/C gnd _4162_/Y vdd OAI21X1
X_4093_ _3873_/A _4098_/S _4101_/C gnd _4094_/A vdd OAI21X1
X_3113_ _3112_/Y _3111_/Y gnd _3113_/Y vdd AND2X2
X_3044_ gnd gnd _3045_/C vdd INVX1
X_2828_ _2828_/A _2776_/Y gnd _2831_/B vdd OR2X2
X_3877_ _3877_/A _3896_/B gnd _3878_/C vdd NOR2X1
X_3946_ _4124_/A _4124_/B _4036_/B gnd _3946_/Y vdd MUX2X1
XSFILL44720x22100 gnd vdd FILL
X_2759_ _2759_/A _2759_/B gnd _2967_/A vdd NAND2X1
X_4429_ _4429_/Q _4431_/CLK _4429_/D gnd vdd DFFPOSX1
XBUFX2_insert8 _3772_/Y gnd _3802_/B vdd BUFX2
X_3800_ _3692_/A _3803_/B _3800_/C gnd _3800_/Y vdd OAI21X1
X_3731_ _3764_/A _3737_/B _3731_/C gnd _4372_/D vdd OAI21X1
X_3662_ _3813_/A _3685_/B _3662_/C gnd _4395_/D vdd AOI21X1
X_2544_ _2331_/A gnd _2544_/Y vdd INVX1
X_3593_ _2986_/B _3616_/B gnd _3593_/Y vdd NAND2X1
X_2613_ _2899_/A gnd _2613_/Y vdd INVX1
X_2475_ _2204_/A _2201_/B gnd _2475_/Y vdd XNOR2X1
X_4076_ _4327_/Q _4012_/S _4010_/C gnd _4077_/A vdd OAI21X1
X_4214_ _4214_/A _4241_/S _4243_/C gnd _4215_/A vdd OAI21X1
XSFILL14480x4100 gnd vdd FILL
X_4145_ _4144_/Y _4145_/B _4155_/C _4142_/Y gnd _4150_/B vdd OAI22X1
X_3027_ gnd gnd _3027_/Y vdd INVX1
X_3929_ _2932_/B _3951_/B _3951_/C gnd _3929_/Y vdd OAI21X1
XFILL70960x12100 gnd vdd FILL
XSFILL14640x16100 gnd vdd FILL
XBUFX2_insert70 _3872_/Y gnd _3904_/B vdd BUFX2
XBUFX2_insert92 _3644_/Q gnd _4036_/B vdd BUFX2
XBUFX2_insert81 _4430_/Q gnd _2361_/B vdd BUFX2
X_2260_ _2255_/Y _2259_/B _2256_/Y gnd _2262_/A vdd AOI21X1
X_2191_ _2191_/A _2191_/B gnd _2191_/Y vdd NAND2X1
XSFILL44240x34100 gnd vdd FILL
XBUFX2_insert291 reset gnd _4206_/C vdd BUFX2
X_3645_ _3645_/Q _4431_/CLK _3570_/Y gnd vdd DFFPOSX1
X_3714_ _3706_/A _3726_/B _3714_/C gnd _3715_/C vdd OAI21X1
XBUFX2_insert280 _3645_/Q gnd _3909_/C vdd BUFX2
X_2527_ _2516_/Y _2519_/Y _2526_/Y gnd _2528_/C vdd OAI21X1
X_2458_ _2451_/C _2458_/B _2458_/C gnd _2539_/B vdd AOI21X1
X_3576_ _3576_/A _3576_/B _3570_/C gnd _3576_/Y vdd AOI21X1
X_4059_ _4059_/A _4057_/Y _4021_/C _4059_/D gnd _4060_/A vdd OAI22X1
X_4128_ _4128_/A _4128_/B _4205_/S gnd _4130_/A vdd MUX2X1
X_2389_ _2429_/A _2429_/B gnd _2391_/A vdd XOR2X1
XSFILL59280x50100 gnd vdd FILL
XCLKBUF1_insert26 clock gnd _4407_/CLK vdd CLKBUF1
XSFILL59760x28100 gnd vdd FILL
X_3292_ _3292_/A _3267_/C _3292_/C gnd _3296_/B vdd NAND3X1
X_3361_ _3360_/Y _3361_/B gnd _3380_/A vdd NOR2X1
X_3430_ _2965_/A _2965_/B gnd _3508_/C vdd AND2X2
X_2312_ _2312_/A _2346_/B gnd _2314_/A vdd NOR2X1
X_2243_ _2242_/Y _2243_/B gnd _2249_/B vdd NOR2X1
XSFILL59440x10100 gnd vdd FILL
X_2174_ _2301_/B _2301_/A gnd _2180_/C vdd AND2X2
XSFILL44720x30100 gnd vdd FILL
X_3628_ _3557_/B _4300_/CLK _3611_/Y gnd vdd DFFPOSX1
X_3559_ _4628_/A _3559_/B gnd _4617_/A vdd AND2X2
XSFILL14160x28100 gnd vdd FILL
X_2861_ _2852_/Y _2860_/Y gnd _2861_/Y vdd NOR2X1
X_2930_ _2930_/A _2920_/Y _2930_/C gnd _2938_/B vdd OAI21X1
X_4600_ _4586_/A _4600_/B gnd _4600_/Y vdd NAND2X1
X_4531_ _4529_/Y _4531_/B _4557_/C gnd _4531_/Y vdd AOI21X1
X_4462_ _4462_/A _4462_/B gnd _4558_/B vdd NOR2X1
X_3413_ _3413_/A _3649_/A gnd _3421_/D vdd AND2X2
X_2792_ _2442_/A _2792_/B gnd _2841_/A vdd NOR2X1
X_2226_ _2226_/A _2226_/B gnd _2227_/B vdd NOR2X1
X_3344_ _3344_/A _3188_/B _3188_/C gnd _3348_/B vdd NAND3X1
X_3275_ _3270_/Y _3275_/B gnd _3275_/Y vdd NOR2X1
X_4393_ _4393_/Q _4298_/CLK _3656_/Y gnd vdd DFFPOSX1
X_2157_ _2140_/A _4250_/A gnd _2157_/Y vdd NAND2X1
XSFILL44560x100 gnd vdd FILL
X_2088_ _2088_/A gnd adrs_bus[2] vdd BUFX2
XFILL70960x20100 gnd vdd FILL
XSFILL14640x24100 gnd vdd FILL
X_3060_ gnd _3372_/B _3372_/C gnd _3061_/A vdd NAND3X1
X_3893_ _4025_/A _3893_/B gnd _3893_/Y vdd NOR2X1
X_2844_ _2789_/Y _2843_/Y _2844_/C _2826_/Y gnd _2844_/Y vdd AOI22X1
X_2913_ _2190_/A _2889_/Y _2913_/C _2913_/D gnd _2913_/Y vdd OAI22X1
X_3962_ _2428_/A _4152_/B _3951_/C gnd _3962_/Y vdd OAI21X1
X_2775_ _2673_/A gnd _2776_/D vdd INVX1
X_4514_ _4493_/C _4499_/Y _4489_/C gnd _4514_/Y vdd NOR3X1
X_4445_ _4445_/Q _4431_/CLK _4445_/D gnd vdd DFFPOSX1
X_4376_ _4376_/Q _4345_/CLK _3807_/Y gnd vdd DFFPOSX1
XSFILL29680x40100 gnd vdd FILL
X_3258_ gnd gnd _3260_/A vdd INVX1
X_3189_ _3189_/A _3345_/B _3188_/B gnd _3191_/B vdd NAND3X1
X_3327_ _3327_/A _3327_/B gnd _3328_/C vdd NOR2X1
X_2209_ _2208_/Y _2207_/Y gnd _2209_/Y vdd NOR2X1
XBUFX2_insert109 _4452_/Q gnd _2856_/A vdd BUFX2
XSFILL59760x36100 gnd vdd FILL
X_4230_ _3799_/A _4389_/Q _4252_/S gnd _4233_/D vdd MUX2X1
X_2560_ _2283_/A _2560_/B gnd _2560_/Y vdd XOR2X1
X_2491_ _2482_/Y _2491_/B _2491_/C gnd _2492_/C vdd AOI21X1
X_3043_ _2342_/Y gnd _3043_/Y vdd INVX1
X_4092_ _3840_/A _4158_/B gnd _4092_/Y vdd NOR2X1
X_4161_ _4161_/A _4161_/B _4205_/S gnd _4163_/A vdd MUX2X1
X_3112_ gnd _3164_/B _3164_/C gnd _3112_/Y vdd NAND3X1
X_3945_ _3945_/A _3943_/Y _3934_/C _3945_/D gnd _3950_/B vdd OAI22X1
X_2827_ _2789_/A gnd _2837_/B vdd INVX1
X_2758_ _2569_/A _2758_/B _2758_/C _2757_/Y gnd _2759_/A vdd AOI22X1
X_3876_ _3843_/A _3879_/B _3875_/Y gnd _3876_/Y vdd AOI21X1
X_4359_ _4359_/Q _4359_/CLK _3804_/Y gnd vdd DFFPOSX1
X_2689_ _2881_/D gnd _2690_/D vdd INVX1
X_4428_ _4428_/Q _4431_/CLK _4428_/D gnd vdd DFFPOSX1
XSFILL59440x8100 gnd vdd FILL
XSFILL14160x36100 gnd vdd FILL
XBUFX2_insert9 _3839_/Y gnd _3846_/B vdd BUFX2
X_3730_ _3726_/A _3726_/B _4042_/A gnd _3731_/C vdd OAI21X1
X_3661_ _4124_/B _3685_/B gnd _3662_/C vdd NOR2X1
X_3592_ _3575_/A data_in[12] gnd _3594_/B vdd NAND2X1
X_2612_ _2706_/B gnd _2612_/Y vdd INVX1
X_2543_ _2533_/Y _2542_/Y _2532_/Y gnd _2549_/A vdd OAI21X1
X_4213_ _3862_/A _4231_/B gnd _4215_/B vdd NOR2X1
X_2474_ _2474_/A _2488_/C _2538_/B _2474_/D gnd _2476_/A vdd AOI22X1
X_4075_ _4253_/A _4020_/B gnd _4075_/Y vdd NOR2X1
X_3026_ _3024_/Y _3130_/B _3026_/C _3130_/D gnd _3030_/A vdd OAI22X1
X_4144_ _3966_/A _4166_/B _4155_/C gnd _4144_/Y vdd OAI21X1
X_3928_ _3928_/A _3928_/B _4027_/S gnd _3930_/A vdd MUX2X1
X_3859_ _4283_/A _3870_/B _3859_/C gnd _4305_/D vdd OAI21X1
XSFILL59280x48100 gnd vdd FILL
XBUFX2_insert60 _4436_/Q gnd _2351_/B vdd BUFX2
XBUFX2_insert71 _3872_/Y gnd _3896_/B vdd BUFX2
XBUFX2_insert82 _4430_/Q gnd _2204_/A vdd BUFX2
XSFILL44560x6100 gnd vdd FILL
XBUFX2_insert93 _3644_/Q gnd _3920_/S vdd BUFX2
X_2190_ _2190_/A _2190_/B gnd _2191_/B vdd OR2X2
XBUFX2_insert281 _3645_/Q gnd _4021_/C vdd BUFX2
XBUFX2_insert292 reset gnd _4239_/C vdd BUFX2
XBUFX2_insert270 _2960_/Y gnd _3345_/B vdd BUFX2
X_3713_ _3813_/A _3737_/B _3712_/Y gnd _3713_/Y vdd OAI21X1
X_3644_ _3644_/Q _4300_/CLK _3567_/Y gnd vdd DFFPOSX1
X_3575_ _3575_/A data_in[5] gnd _3576_/B vdd NAND2X1
X_2526_ _2520_/Y gnd _2526_/Y vdd INVX1
X_2388_ _2388_/A _2388_/B gnd _2400_/A vdd NOR2X1
X_2457_ _2456_/A _2455_/Y gnd _2458_/C vdd NOR2X1
X_4058_ _4341_/Q _4074_/S _4021_/C gnd _4059_/A vdd OAI21X1
X_4127_ _4126_/Y _4127_/B _4247_/C _4124_/Y gnd _4128_/A vdd OAI22X1
XSFILL44720x28100 gnd vdd FILL
X_3009_ _3009_/A _3007_/Y gnd _3010_/C vdd AND2X2
XSFILL44400x10100 gnd vdd FILL
XSFILL14320x4100 gnd vdd FILL
XCLKBUF1_insert27 clock gnd _4300_/CLK vdd CLKBUF1
XFILL71120x12100 gnd vdd FILL
X_2242_ _2252_/A _2252_/B gnd _2242_/Y vdd NOR2X1
X_3291_ gnd _3343_/B gnd _3291_/Y vdd NAND2X1
X_3360_ _3360_/A _3204_/B _3359_/Y _3204_/D gnd _3360_/Y vdd OAI22X1
X_2311_ _2311_/A _2310_/Y gnd _2311_/Y vdd NOR2X1
X_2173_ _2168_/Y _2172_/B _2171_/B gnd _2177_/A vdd AOI21X1
X_2509_ _2497_/Y _2505_/Y gnd _2509_/Y vdd NAND2X1
X_3627_ _3556_/B _3632_/CLK _3609_/Y gnd vdd DFFPOSX1
X_3558_ _4628_/A _3545_/A gnd _4614_/A vdd AND2X2
X_3489_ _3483_/Y _3488_/Y gnd _3489_/Y vdd NAND2X1
X_2860_ _2857_/Y _2859_/Y _2855_/Y gnd _2860_/Y vdd NAND3X1
X_2791_ _2442_/A _2792_/B gnd _2795_/C vdd NAND2X1
X_4530_ _4558_/B _4530_/B _4575_/Q _4556_/D gnd _4531_/B vdd AOI22X1
X_4461_ _4560_/A gnd _4462_/B vdd INVX1
X_3412_ _3402_/Y _3417_/D gnd _3419_/D vdd NOR2X1
X_4392_ _4392_/Q _4394_/CLK _3653_/Y gnd vdd DFFPOSX1
X_2225_ _2228_/A _2786_/A gnd _2226_/A vdd NOR2X1
X_3343_ gnd _3343_/B gnd _3348_/A vdd NAND2X1
X_3274_ _3272_/Y _3274_/B _3273_/Y gnd _3275_/B vdd NAND3X1
X_2087_ _2161_/Y gnd adrs_bus[15] vdd BUFX2
X_2156_ _4556_/C gnd _2158_/B vdd INVX1
XSFILL29680x38100 gnd vdd FILL
X_2989_ _2980_/Y _2989_/B gnd _2990_/C vdd NOR2X1
XSFILL29360x20100 gnd vdd FILL
XSFILL14640x40100 gnd vdd FILL
X_2912_ _2907_/Y _2901_/Y _2912_/C gnd _2912_/Y vdd OAI21X1
X_3961_ _3961_/A _3961_/B _4027_/S gnd _3963_/A vdd MUX2X1
X_2774_ _2829_/B gnd _2776_/B vdd INVX1
X_3892_ _4283_/A _3893_/B _3892_/C gnd _3892_/Y vdd AOI21X1
X_4513_ _4506_/C _4513_/B _4513_/C gnd _4516_/B vdd OAI21X1
X_2843_ _2838_/Y _2825_/A _2842_/Y gnd _2843_/Y vdd NOR3X1
XSFILL59440x16100 gnd vdd FILL
X_4375_ _4253_/A _4359_/CLK _4375_/D gnd vdd DFFPOSX1
X_3326_ _3324_/Y _3326_/B _3325_/Y gnd _3327_/B vdd NAND3X1
X_4444_ _4444_/Q _4431_/CLK _4444_/D gnd vdd DFFPOSX1
X_2139_ _2140_/A _4184_/A gnd _2139_/Y vdd NAND2X1
XSFILL44720x36100 gnd vdd FILL
X_3257_ _3256_/Y _3257_/B gnd _3276_/A vdd NOR2X1
X_3188_ _3188_/A _3188_/B _3188_/C gnd _3192_/B vdd NAND3X1
X_2208_ _2346_/B _2312_/A gnd _2208_/Y vdd NOR2X1
XSFILL59760x52100 gnd vdd FILL
X_2490_ _2482_/B _2490_/B gnd _2491_/C vdd NOR2X1
X_4160_ _4159_/Y _4158_/Y _4101_/C _4160_/D gnd _4161_/A vdd OAI22X1
XFILL71120x20100 gnd vdd FILL
X_3111_ _2192_/Y _2977_/B _3090_/B gnd _3111_/Y vdd NAND3X1
X_4091_ _4408_/Q _4392_/Q _4098_/S gnd _4094_/D vdd MUX2X1
X_3042_ _3023_/Y _3042_/B _3041_/Y gnd _3042_/Y vdd NAND3X1
X_3944_ _3944_/A _4030_/S _3909_/C gnd _3945_/A vdd OAI21X1
X_3875_ _4329_/Q _3879_/B gnd _3875_/Y vdd NOR2X1
X_2826_ _2789_/Y _2825_/Y gnd _2826_/Y vdd NAND2X1
X_2688_ _2693_/B gnd _2690_/A vdd INVX1
X_2757_ _2703_/A _2703_/B _2756_/Y gnd _2757_/Y vdd NOR3X1
X_4358_ _4241_/A _4407_/CLK _3802_/Y gnd vdd DFFPOSX1
X_4289_ _3764_/A _4287_/B _4288_/Y gnd _4289_/Y vdd AOI21X1
X_3309_ _3309_/A _3309_/B gnd _3328_/A vdd NOR2X1
XSFILL59920x12100 gnd vdd FILL
X_4427_ _4427_/Q _4297_/CLK _4427_/D gnd vdd DFFPOSX1
XSFILL14160x52100 gnd vdd FILL
X_2542_ _2558_/A _2528_/Y gnd _2542_/Y vdd AND2X2
X_3591_ _3591_/A _3589_/Y _3579_/C gnd _3591_/Y vdd AOI21X1
X_2611_ _2609_/Y _2301_/A _2611_/C _2899_/A gnd _2615_/A vdd AOI22X1
X_3660_ _3454_/Y gnd _3813_/A vdd INVX4
X_4212_ _4212_/A _4212_/B _4241_/S gnd _4212_/Y vdd MUX2X1
X_2473_ _2461_/B _2473_/B gnd _2538_/B vdd NOR2X1
X_4143_ _4365_/Q _4088_/B gnd _4145_/B vdd NOR2X1
XSFILL14320x12100 gnd vdd FILL
X_4074_ _4359_/Q _3836_/A _4074_/S gnd _4077_/D vdd MUX2X1
X_3025_ gnd gnd _3026_/C vdd INVX1
X_3858_ _4191_/A _3870_/B gnd _3859_/C vdd NAND2X1
X_3927_ _3927_/A _3925_/Y _3934_/C _3927_/D gnd _3928_/A vdd OAI22X1
XSFILL29680x46100 gnd vdd FILL
X_3789_ _4352_/Q _3792_/B gnd _3789_/Y vdd NAND2X1
XSFILL30160x34100 gnd vdd FILL
X_2809_ _2201_/B gnd _2810_/D vdd INVX1
XBUFX2_insert61 _4436_/Q gnd _2768_/A vdd BUFX2
XBUFX2_insert50 _3805_/Y gnd _3832_/B vdd BUFX2
XBUFX2_insert72 _4442_/Q gnd _2104_/A vdd BUFX2
XBUFX2_insert83 _4430_/Q gnd _4600_/B vdd BUFX2
XBUFX2_insert94 _4427_/Q gnd _2609_/A vdd BUFX2
X_3712_ _3703_/B _3726_/B _4363_/Q gnd _3712_/Y vdd OAI21X1
XBUFX2_insert260 _4440_/Q gnd _2429_/A vdd BUFX2
XBUFX2_insert282 _3645_/Q gnd _4010_/C vdd BUFX2
X_2525_ _2525_/A gnd _2528_/A vdd INVX1
XBUFX2_insert271 _2960_/Y gnd _2961_/A vdd BUFX2
XSFILL59440x24100 gnd vdd FILL
X_3643_ _4085_/A _4300_/CLK _3582_/Y gnd vdd DFFPOSX1
X_3574_ _4166_/B _3574_/B gnd _3576_/A vdd NAND2X1
XBUFX2_insert293 reset gnd _4228_/C vdd BUFX2
X_2387_ _4072_/A _4250_/A gnd _2388_/B vdd XOR2X1
X_4126_ _3948_/A _4124_/S _4111_/C gnd _4126_/Y vdd OAI21X1
X_2456_ _2456_/A _2455_/Y gnd _2458_/B vdd NAND2X1
X_4057_ _4057_/A _4002_/B gnd _4057_/Y vdd NOR2X1
X_3008_ gnd _3372_/B _3372_/C gnd _3009_/A vdd NAND3X1
XCLKBUF1_insert28 clock gnd _4394_/CLK vdd CLKBUF1
X_2241_ _2253_/A _2253_/B gnd _2243_/B vdd NOR2X1
X_3290_ _3290_/A _3289_/Y gnd _3290_/Y vdd NOR2X1
X_2172_ _2168_/Y _2172_/B gnd _2172_/Y vdd XOR2X1
X_2310_ _2361_/A _2361_/B gnd _2310_/Y vdd AND2X2
X_2508_ _2507_/Y gnd _2508_/Y vdd INVX1
X_3488_ _3495_/A _3487_/Y _3485_/Y gnd _3488_/Y vdd NAND3X1
X_3626_ _3555_/A _3632_/CLK _3626_/D gnd vdd DFFPOSX1
X_3557_ _3561_/A _3557_/B gnd _4611_/A vdd AND2X2
X_4109_ _4109_/A _4378_/Q _4124_/S gnd _4112_/D vdd MUX2X1
X_2439_ _2442_/A _2442_/B gnd _2443_/B vdd NAND2X1
XSFILL44400x6100 gnd vdd FILL
XSFILL59920x20100 gnd vdd FILL
XSFILL29360x18100 gnd vdd FILL
X_2790_ _2906_/A gnd _2792_/B vdd INVX1
X_4391_ _3836_/A _4359_/CLK _4391_/D gnd vdd DFFPOSX1
X_3342_ _3338_/Y _3342_/B gnd _3354_/B vdd NOR2X1
X_4460_ _4460_/A _4548_/C gnd _4460_/Y vdd NAND2X1
X_3411_ _3401_/C gnd _3649_/C vdd INVX1
XSFILL14320x20100 gnd vdd FILL
X_2224_ _2222_/Y _2223_/Y gnd _2226_/B vdd NOR2X1
X_2155_ _2151_/A _2153_/Y _2155_/C gnd _2155_/Y vdd OAI21X1
X_3273_ _3143_/A gnd gnd _3143_/D gnd _3273_/Y vdd AOI22X1
X_2086_ _2158_/Y gnd adrs_bus[14] vdd BUFX2
X_2988_ _2988_/A _2983_/Y _2988_/C gnd _2989_/B vdd NAND3X1
X_3609_ _3609_/A _3607_/Y _3615_/C gnd _3609_/Y vdd AOI21X1
X_4589_ _4594_/A _4589_/B _4588_/Y gnd _4589_/Y vdd OAI21X1
XSFILL44400x16100 gnd vdd FILL
XFILL71120x18100 gnd vdd FILL
X_3891_ _4337_/Q _3893_/B gnd _3892_/C vdd NOR2X1
X_3960_ _3960_/A _3960_/B _3982_/C _3960_/D gnd _3961_/A vdd OAI22X1
X_2911_ _2909_/Y _2910_/Y _2911_/C gnd _2912_/C vdd AOI21X1
X_2773_ _2769_/Y _2773_/B _2766_/Y gnd _2789_/A vdd NAND3X1
X_4512_ _2138_/A gnd _4513_/C vdd INVX1
X_2842_ _2842_/A _2619_/A _2841_/Y gnd _2842_/Y vdd OAI21X1
X_4374_ _4064_/A _4407_/CLK _3735_/Y gnd vdd DFFPOSX1
X_3256_ _3256_/A _3204_/B _3256_/C _3204_/D gnd _3256_/Y vdd OAI22X1
XSFILL59440x32100 gnd vdd FILL
X_3325_ _3143_/A gnd gnd _3143_/D gnd _3325_/Y vdd AOI22X1
X_4443_ _4443_/Q _4431_/CLK _4443_/D gnd vdd DFFPOSX1
X_2138_ _2138_/A gnd _2138_/Y vdd INVX1
X_3187_ gnd _3343_/B gnd _3187_/Y vdd NAND2X1
X_2207_ _2346_/B _2312_/A gnd _2207_/Y vdd AND2X2
XSFILL44720x52100 gnd vdd FILL
X_3110_ _2308_/Y _3194_/B _3110_/C gnd _3110_/Y vdd NAND3X1
X_4090_ _4090_/A _4090_/B _4155_/C _4090_/D gnd _4095_/B vdd OAI22X1
X_3041_ _3036_/Y _3041_/B gnd _3041_/Y vdd NOR2X1
X_3943_ _4363_/Q _3943_/B gnd _3943_/Y vdd NOR2X1
X_2825_ _2825_/A _2807_/Y _2825_/C gnd _2825_/Y vdd OAI21X1
X_3874_ _3740_/A _3879_/B _3873_/Y gnd _4328_/D vdd AOI21X1
X_2687_ _2671_/Y _2687_/B gnd _2744_/A vdd NAND2X1
X_2756_ _2706_/Y _2756_/B _2755_/Y gnd _2756_/Y vdd NAND3X1
X_4426_ _4426_/Q _4297_/CLK _4426_/D gnd vdd DFFPOSX1
X_4357_ _3799_/A _4407_/CLK _3800_/Y gnd vdd DFFPOSX1
X_3239_ gnd _3343_/B gnd _3244_/A vdd NAND2X1
X_3308_ _3308_/A _3204_/B _3307_/Y _3204_/D gnd _3309_/A vdd OAI22X1
X_4288_ _4045_/A _4287_/B gnd _4288_/Y vdd NOR2X1
X_3590_ _3699_/A _3590_/B gnd _3591_/A vdd NAND2X1
X_2472_ _2465_/A _2465_/B _2472_/C gnd _2488_/C vdd OAI21X1
X_2541_ _2541_/A _2539_/Y _2541_/C gnd _2558_/A vdd OAI21X1
X_2610_ _2298_/B gnd _2611_/C vdd INVX1
X_4073_ _4071_/Y _4040_/B _4072_/Y gnd _4073_/Y vdd AOI21X1
X_4211_ _4210_/Y _4209_/Y _4243_/C _4211_/D gnd _4211_/Y vdd OAI22X1
X_4142_ _4142_/A _3816_/A _4153_/S gnd _4142_/Y vdd MUX2X1
X_3024_ gnd gnd _3024_/Y vdd INVX1
X_3857_ _4281_/A _3862_/B _3856_/Y gnd _4304_/D vdd OAI21X1
X_2808_ _2482_/B gnd _2822_/B vdd INVX1
X_3788_ _3788_/A _3775_/B _3787_/Y gnd _3788_/Y vdd OAI21X1
X_3926_ _4329_/Q _3992_/B _3934_/C gnd _3927_/A vdd OAI21X1
X_2739_ _2660_/Y _4072_/A _2739_/C _2737_/Y gnd _2748_/A vdd AOI22X1
X_4409_ _4266_/A _4394_/CLK _4267_/Y gnd vdd DFFPOSX1
XSFILL44400x24100 gnd vdd FILL
XSFILL28880x14100 gnd vdd FILL
XBUFX2_insert40 _3738_/Y gnd _3767_/B vdd BUFX2
XBUFX2_insert62 _4436_/Q gnd _4228_/A vdd BUFX2
XBUFX2_insert51 _3805_/Y gnd _3823_/B vdd BUFX2
XBUFX2_insert84 _4430_/Q gnd _2880_/A vdd BUFX2
XBUFX2_insert73 _4442_/Q gnd _2899_/A vdd BUFX2
XBUFX2_insert95 _4427_/Q gnd _2301_/B vdd BUFX2
XSFILL60240x46100 gnd vdd FILL
XBUFX2_insert283 _3645_/Q gnd _4065_/C vdd BUFX2
X_3711_ _3811_/A _3737_/B _3710_/Y gnd _3711_/Y vdd OAI21X1
X_3642_ _3642_/Q _4300_/CLK _3579_/Y gnd vdd DFFPOSX1
XBUFX2_insert261 _4440_/Q gnd _2794_/A vdd BUFX2
XBUFX2_insert250 _4443_/Q gnd _2377_/A vdd BUFX2
XBUFX2_insert294 reset gnd _3951_/C vdd BUFX2
XBUFX2_insert272 _2960_/Y gnd _3007_/B vdd BUFX2
X_2524_ _2509_/Y _2525_/A gnd _2529_/A vdd OR2X2
X_2455_ _2799_/A gnd _2455_/Y vdd INVX1
X_3573_ _3573_/A _3573_/B _3582_/C gnd _3646_/D vdd AOI21X1
X_4056_ _4056_/A _3691_/A _4074_/S gnd _4059_/D vdd MUX2X1
X_2386_ _2848_/A _4261_/A gnd _2388_/A vdd XOR2X1
X_4125_ _3947_/A _4180_/B gnd _4127_/B vdd NOR2X1
X_3007_ _2167_/Y _3007_/B _3032_/B gnd _3007_/Y vdd NAND3X1
X_3909_ _4312_/Q _3920_/S _3909_/C gnd _3909_/Y vdd OAI21X1
XSFILL59920x18100 gnd vdd FILL
XSFILL43920x12100 gnd vdd FILL
XCLKBUF1_insert29 clock gnd _4431_/CLK vdd CLKBUF1
X_2240_ _2252_/B gnd _2253_/B vdd INVX1
X_2171_ _2170_/Y _2171_/B gnd _2172_/B vdd NOR2X1
XSFILL14320x18100 gnd vdd FILL
X_3625_ _3625_/Q _4431_/CLK _3624_/Y gnd vdd DFFPOSX1
X_2507_ _2502_/Y _2496_/Y _2503_/Y gnd _2507_/Y vdd OAI21X1
X_2438_ _2906_/A gnd _2442_/B vdd INVX1
X_3487_ _3487_/A _3508_/B _3508_/C gnd _3487_/Y vdd NAND3X1
X_3556_ _4628_/A _3556_/B gnd _3490_/B vdd AND2X2
X_4039_ _4039_/A _4040_/B _4206_/C gnd _4039_/Y vdd OAI21X1
X_2369_ _2661_/A _2571_/B gnd _3349_/A vdd AND2X2
X_4108_ _4108_/A _4130_/B _4107_/Y gnd _4425_/D vdd AOI21X1
XFILL70960x50100 gnd vdd FILL
X_4390_ _4390_/Q _4407_/CLK _3835_/Y gnd vdd DFFPOSX1
X_3341_ _3341_/A _3341_/B _3341_/C gnd _3342_/B vdd OAI21X1
X_3272_ gnd _3188_/B _3194_/C gnd _3272_/Y vdd NAND3X1
X_3410_ _3410_/A _3410_/B gnd _3410_/Y vdd NOR2X1
X_2085_ _2155_/Y gnd adrs_bus[13] vdd BUFX2
X_2223_ _2830_/B gnd _2223_/Y vdd INVX1
X_2154_ _2151_/A _4239_/A gnd _2155_/C vdd NAND2X1
X_2987_ _3143_/A _2987_/B gnd _3143_/D gnd _2988_/C vdd AOI22X1
X_3608_ _3556_/B _3605_/B gnd _3609_/A vdd NAND2X1
XSFILL14800x14100 gnd vdd FILL
X_4588_ _4594_/A _4588_/B gnd _4588_/Y vdd NAND2X1
X_3539_ _3555_/A gnd _3540_/B vdd INVX1
XSFILL29680x2100 gnd vdd FILL
XSFILL44400x32100 gnd vdd FILL
XSFILL29840x30100 gnd vdd FILL
XFILL71120x34100 gnd vdd FILL
X_3890_ _4281_/A _3896_/B _3889_/Y gnd _4336_/D vdd AOI21X1
X_2841_ _2841_/A _2840_/Y gnd _2841_/Y vdd NOR2X1
X_2910_ _2895_/A _2898_/Y gnd _2910_/Y vdd NAND2X1
X_2772_ _2770_/Y _2772_/B _2772_/C _2768_/A gnd _2773_/B vdd AOI22X1
X_4511_ _4511_/A _4511_/B _4557_/C gnd _4511_/Y vdd AOI21X1
X_4442_ _4442_/Q _4297_/CLK _4442_/D gnd vdd DFFPOSX1
X_4373_ _4231_/A _4373_/CLK _3733_/Y gnd vdd DFFPOSX1
X_3255_ gnd gnd _3256_/C vdd INVX1
X_3324_ gnd _3240_/B _3324_/C gnd _3324_/Y vdd NAND3X1
X_2206_ _2202_/A _2206_/B _2213_/B gnd _2206_/Y vdd AOI21X1
X_2137_ _2140_/A _2137_/B _2136_/Y gnd _2137_/Y vdd OAI21X1
X_3186_ _3182_/Y _3186_/B gnd _3198_/B vdd NOR2X1
XSFILL59920x26100 gnd vdd FILL
X_3040_ _3040_/A _3037_/Y _3040_/C gnd _3041_/B vdd NAND3X1
X_3942_ _4347_/Q _4379_/Q _4030_/S gnd _3945_/D vdd MUX2X1
XSFILL14320x26100 gnd vdd FILL
X_2824_ _2810_/Y _2824_/B _2823_/Y _2814_/Y gnd _2825_/C vdd AOI22X1
X_3873_ _3873_/A _3873_/B gnd _3873_/Y vdd NOR2X1
X_2686_ _2678_/Y _2685_/Y gnd _2687_/B vdd AND2X2
X_4356_ _4041_/A _4298_/CLK _4356_/D gnd vdd DFFPOSX1
X_2755_ _2751_/Y _2752_/Y _2755_/C _2755_/D gnd _2755_/Y vdd AOI22X1
X_4425_ _4425_/Q _4297_/CLK _4425_/D gnd vdd DFFPOSX1
X_4287_ _3729_/A _4287_/B _4286_/Y gnd _4419_/D vdd AOI21X1
X_3307_ gnd gnd _3307_/Y vdd INVX1
X_3238_ _3238_/A _3237_/Y gnd _3250_/B vdd NOR2X1
X_3169_ _3143_/A gnd gnd _3143_/D gnd _3169_/Y vdd AOI22X1
XSFILL29360x42100 gnd vdd FILL
X_2540_ _2525_/A _2509_/Y gnd _2541_/C vdd NOR2X1
X_4210_ _4032_/A _4241_/S _4243_/C gnd _4210_/Y vdd OAI21X1
X_2471_ _2465_/Y _2473_/B gnd _2471_/Y vdd XNOR2X1
X_4072_ _4072_/A _4217_/B _4239_/C gnd _4072_/Y vdd OAI21X1
X_4141_ _4141_/A _4152_/B _4140_/Y gnd _4428_/D vdd AOI21X1
X_3023_ _3022_/Y _3023_/B gnd _3023_/Y vdd NOR2X1
XSFILL59440x38100 gnd vdd FILL
X_3925_ _4297_/Q _3943_/B gnd _3925_/Y vdd NOR2X1
X_2738_ _2848_/A _4261_/A gnd _2739_/C vdd NAND2X1
X_3856_ _4002_/A _3862_/B gnd _3856_/Y vdd NAND2X1
X_2807_ _2838_/A _2795_/Y _2806_/Y gnd _2807_/Y vdd AOI21X1
X_3787_ _4351_/Q _3775_/B gnd _3787_/Y vdd NAND2X1
X_2669_ _4228_/A _2669_/B gnd _2669_/Y vdd NAND2X1
X_4339_ _4214_/A _4373_/CLK _3896_/Y gnd vdd DFFPOSX1
XSFILL14800x22100 gnd vdd FILL
X_4408_ _4408_/Q _4345_/CLK _4265_/Y gnd vdd DFFPOSX1
XSFILL44400x40100 gnd vdd FILL
XBUFX2_insert41 _4448_/Q gnd _2218_/B vdd BUFX2
XBUFX2_insert63 _2968_/Y gnd _3346_/B vdd BUFX2
XBUFX2_insert85 _4430_/Q gnd _2916_/A vdd BUFX2
XBUFX2_insert96 _4427_/Q gnd _2799_/A vdd BUFX2
XSFILL13840x100 gnd vdd FILL
XBUFX2_insert74 _4442_/Q gnd _2406_/A vdd BUFX2
XBUFX2_insert52 _3805_/Y gnd _3809_/B vdd BUFX2
XBUFX2_insert251 _4434_/Q gnd _4206_/A vdd BUFX2
X_3710_ _3703_/B _3726_/B _3932_/A gnd _3710_/Y vdd OAI21X1
X_3572_ _3575_/A data_in[4] gnd _3573_/B vdd NAND2X1
XBUFX2_insert262 _4440_/Q gnd _2713_/A vdd BUFX2
XBUFX2_insert240 _4446_/Q gnd _2881_/D vdd BUFX2
XBUFX2_insert295 reset gnd _3649_/A vdd BUFX2
X_3641_ _3641_/Q _4297_/CLK _3576_/Y gnd vdd DFFPOSX1
XBUFX2_insert284 _3645_/Q gnd _3982_/C vdd BUFX2
XBUFX2_insert273 _4087_/Y gnd _4158_/B vdd BUFX2
X_2523_ _2511_/Y _2522_/B gnd _2525_/A vdd NAND2X1
X_2385_ _2373_/Y _2385_/B _2384_/Y gnd _2385_/Y vdd NAND3X1
X_2454_ _2445_/B _2452_/Y gnd _2459_/B vdd NAND2X1
X_4055_ _4055_/A _4053_/Y _4021_/C _4055_/D gnd _4055_/Y vdd OAI22X1
X_4124_ _4124_/A _4124_/B _4124_/S gnd _4124_/Y vdd MUX2X1
X_3006_ _3006_/A _3032_/B _2947_/A gnd _3006_/Y vdd NAND3X1
X_3908_ _4360_/Q _3921_/B gnd _3910_/B vdd NOR2X1
X_3839_ _3839_/A _3703_/Y gnd _3839_/Y vdd NAND2X1
XSFILL60400x22100 gnd vdd FILL
X_2170_ _2298_/B _2298_/A gnd _2170_/Y vdd NOR2X1
XSFILL29040x14100 gnd vdd FILL
XSFILL14320x34100 gnd vdd FILL
X_3624_ _3623_/Y _3624_/B _3570_/C gnd _3624_/Y vdd AOI21X1
X_3555_ _3555_/A _3561_/A gnd _4605_/A vdd AND2X2
X_2506_ _2500_/Y _2505_/Y gnd _3202_/A vdd XOR2X1
X_2368_ _2331_/A _2330_/B gnd _3323_/A vdd AND2X2
X_2437_ _2906_/A _2437_/B gnd _2440_/A vdd NAND2X1
X_3486_ data_in[8] gnd _3487_/A vdd INVX1
X_4038_ _4037_/Y _4038_/B _4027_/S gnd _4038_/Y vdd MUX2X1
X_4107_ _4585_/B _4130_/B _4162_/C gnd _4107_/Y vdd OAI21X1
X_2299_ _2297_/Y _2298_/Y gnd _2299_/Y vdd NOR2X1
XSFILL29360x50100 gnd vdd FILL
XSFILL29840x28100 gnd vdd FILL
X_2222_ _2228_/A gnd _2222_/Y vdd INVX1
X_3271_ _3271_/A _3141_/B gnd _3274_/B vdd NAND2X1
X_3340_ gnd _3340_/B gnd _3341_/C vdd NAND2X1
X_2084_ _2152_/Y gnd adrs_bus[12] vdd BUFX2
X_2153_ _4578_/Q gnd _2153_/Y vdd INVX1
XSFILL29520x10100 gnd vdd FILL
X_2986_ _2986_/A _2986_/B _2986_/C gnd _3143_/A vdd NOR3X1
XSFILL14800x30100 gnd vdd FILL
X_3607_ _3601_/A data_in[1] gnd _3607_/Y vdd NAND2X1
X_3538_ _3538_/A _3537_/Y gnd _3538_/Y vdd NAND2X1
X_4587_ _3441_/B gnd _4589_/B vdd INVX1
X_3469_ _3422_/B _3469_/B gnd _3469_/Y vdd NAND2X1
XFILL71120x50100 gnd vdd FILL
X_2771_ _2100_/A gnd _2772_/C vdd INVX1
X_2840_ _2794_/A _2794_/B _2795_/C gnd _2840_/Y vdd OAI21X1
X_4372_ _4042_/A _4436_/CLK _4372_/D gnd vdd DFFPOSX1
X_4510_ _4558_/B _4604_/Y _2135_/A _4556_/D gnd _4511_/B vdd AOI22X1
X_4441_ _4441_/Q _4431_/CLK _4441_/D gnd vdd DFFPOSX1
X_3254_ _2522_/Y gnd _3256_/A vdd INVX1
XSFILL58960x34100 gnd vdd FILL
X_3323_ _3323_/A _3141_/B gnd _3326_/B vdd NAND2X1
X_3185_ _3185_/A _3341_/B _3184_/Y gnd _3186_/B vdd OAI21X1
X_2205_ _2204_/Y _2213_/B gnd _2206_/B vdd NOR2X1
X_2136_ _2124_/A _2136_/B gnd _2136_/Y vdd NAND2X1
X_2969_ _3294_/B _2969_/B gnd _3341_/B vdd NAND2X1
XSFILL45200x8100 gnd vdd FILL
X_3941_ _3941_/A _3941_/B _3940_/Y gnd _4442_/D vdd AOI21X1
XSFILL29520x2100 gnd vdd FILL
X_2823_ _2823_/A _2817_/Y gnd _2823_/Y vdd NOR2X1
X_2754_ _2292_/B _2290_/B gnd _2755_/D vdd NAND2X1
X_3872_ _3651_/A _3839_/A gnd _3872_/Y vdd AND2X2
X_2685_ _2735_/C _2684_/Y gnd _2685_/Y vdd NOR2X1
X_3306_ _3306_/A gnd _3308_/A vdd INVX1
X_4355_ _4208_/A _4373_/CLK _3796_/Y gnd vdd DFFPOSX1
XSFILL60080x2100 gnd vdd FILL
X_4424_ _4424_/Q _4431_/CLK _4424_/D gnd vdd DFFPOSX1
X_4286_ _4212_/A _4287_/B gnd _4286_/Y vdd NOR2X1
X_3237_ _3235_/Y _3341_/B _3237_/C gnd _3237_/Y vdd OAI21X1
X_2119_ _2118_/A _2119_/B _2119_/C gnd _2081_/A vdd OAI21X1
X_3168_ gnd _3194_/B _3116_/C gnd _3168_/Y vdd NAND3X1
X_3099_ gnd gnd _3100_/C vdd INVX1
XSFILL29680x8100 gnd vdd FILL
XSFILL29840x36100 gnd vdd FILL
X_2470_ _2474_/A _2472_/C gnd _2473_/B vdd NAND2X1
X_4140_ _2127_/B _4152_/B _3951_/C gnd _4140_/Y vdd OAI21X1
X_4071_ _4071_/A _4071_/B _4027_/S gnd _4071_/Y vdd MUX2X1
X_3022_ _3020_/Y _3204_/B _3022_/C _3204_/D gnd _3022_/Y vdd OAI22X1
X_3924_ _4266_/A _4393_/Q _3992_/B gnd _3927_/D vdd MUX2X1
X_2668_ _2762_/C _2668_/B gnd _2670_/B vdd NAND2X1
X_2737_ _2659_/B _2758_/B gnd _2737_/Y vdd NAND2X1
X_2806_ _2806_/A _2805_/Y _2803_/Y gnd _2806_/Y vdd OAI21X1
X_3855_ _3788_/A _3852_/B _3854_/Y gnd _4303_/D vdd OAI21X1
X_3786_ _3752_/A _3786_/B _3785_/Y gnd _3786_/Y vdd OAI21X1
X_4407_ _4407_/Q _4407_/CLK _3698_/Y gnd vdd DFFPOSX1
X_4338_ _4025_/A _4417_/CLK _4338_/D gnd vdd DFFPOSX1
X_4269_ _3811_/A _4269_/B _4268_/Y gnd _4269_/Y vdd AOI21X1
XSFILL59280x100 gnd vdd FILL
X_2599_ _2599_/A _2915_/A _2916_/A _2599_/D gnd _2600_/B vdd AOI22X1
XBUFX2_insert42 _4448_/Q gnd _2421_/A vdd BUFX2
XBUFX2_insert20 _3564_/Y gnd _3574_/B vdd BUFX2
XBUFX2_insert53 _3805_/Y gnd _3819_/B vdd BUFX2
XBUFX2_insert86 _3644_/Q gnd _3968_/S vdd BUFX2
XBUFX2_insert75 _4442_/Q gnd _2298_/A vdd BUFX2
XSFILL59600x14100 gnd vdd FILL
XBUFX2_insert97 _4427_/Q gnd _4591_/B vdd BUFX2
XBUFX2_insert64 _2968_/Y gnd _3372_/B vdd BUFX2
XBUFX2_insert252 _4434_/Q gnd _2778_/A vdd BUFX2
XBUFX2_insert230 _4449_/Q gnd _2830_/B vdd BUFX2
X_2522_ _2517_/Y _2522_/B gnd _2522_/Y vdd XOR2X1
XBUFX2_insert285 _3645_/Q gnd _4004_/C vdd BUFX2
X_3640_ _3699_/A _4300_/CLK _3591_/Y gnd vdd DFFPOSX1
X_3571_ _3905_/A _3590_/B gnd _3573_/A vdd NAND2X1
XBUFX2_insert241 _4446_/Q gnd _2418_/A vdd BUFX2
XBUFX2_insert263 _4440_/Q gnd _2290_/B vdd BUFX2
XBUFX2_insert296 reset gnd _4162_/C vdd BUFX2
XBUFX2_insert274 _4087_/Y gnd _4088_/B vdd BUFX2
X_4123_ _4123_/A _4123_/B _4111_/C _4123_/D gnd _4128_/B vdd OAI22X1
X_2384_ _2377_/Y _2378_/Y _2384_/C gnd _2384_/Y vdd NOR3X1
X_2453_ _2451_/Y _2452_/Y gnd _2453_/Y vdd XNOR2X1
X_4054_ _4232_/A _4052_/S _4065_/C gnd _4055_/A vdd OAI21X1
X_3005_ gnd _3343_/B gnd _3005_/Y vdd NAND2X1
X_3907_ _4030_/S gnd _3907_/Y vdd INVX8
X_3838_ _3699_/A _3700_/Y gnd _3839_/A vdd NOR2X1
X_3769_ _4327_/Q _3760_/B gnd _3770_/C vdd NAND2X1
XSFILL29360x48100 gnd vdd FILL
XSFILL14320x50100 gnd vdd FILL
X_2505_ _2502_/Y _2504_/Y gnd _2505_/Y vdd NOR2X1
X_3485_ _3513_/A _3513_/B _3485_/C gnd _3485_/Y vdd OAI21X1
X_3623_ _3562_/A _3616_/B gnd _3623_/Y vdd NAND2X1
X_3554_ _3561_/A _3554_/B gnd _4602_/A vdd NOR2X1
X_2367_ _2351_/A _2351_/B gnd _3297_/A vdd AND2X2
X_2436_ _2442_/A gnd _2437_/B vdd INVX1
X_2298_ _2298_/A _2298_/B gnd _2298_/Y vdd AND2X2
X_4106_ _4105_/Y _4106_/B _4205_/S gnd _4108_/A vdd MUX2X1
X_4037_ _4036_/Y _4037_/B _4004_/C _4034_/Y gnd _4037_/Y vdd OAI22X1
XFILL71120x48100 gnd vdd FILL
X_2221_ _2218_/Y _2221_/B _2216_/Y gnd _2227_/A vdd OAI21X1
X_2152_ _2151_/A _2152_/B _2151_/Y gnd _2152_/Y vdd OAI21X1
X_3270_ _3270_/A _3270_/B _3269_/Y gnd _3270_/Y vdd NAND3X1
X_2083_ _2149_/Y gnd adrs_bus[11] vdd BUFX2
X_2985_ _2965_/B _2941_/Y _2982_/A gnd _3143_/D vdd NOR3X1
X_3606_ _3606_/A _3606_/B _3615_/C gnd _3626_/D vdd AOI21X1
X_3468_ _3468_/A _3467_/Y gnd _3666_/A vdd NAND2X1
X_4586_ _4586_/A _4586_/B _4585_/Y gnd _4586_/Y vdd OAI21X1
X_3537_ _3495_/A _3536_/Y _3537_/C gnd _3537_/Y vdd NAND3X1
X_3399_ _2986_/B _2986_/A gnd _3410_/A vdd NAND2X1
XSFILL44880x18100 gnd vdd FILL
X_2419_ _2417_/Y _2418_/Y gnd _2419_/Y vdd NAND2X1
X_2770_ _2101_/A gnd _2770_/Y vdd INVX1
X_3322_ _3317_/Y _3322_/B _3321_/Y gnd _3327_/A vdd NAND3X1
X_4371_ _4031_/A _4407_/CLK _4371_/D gnd vdd DFFPOSX1
X_4440_ _4440_/Q _4297_/CLK _4440_/D gnd vdd DFFPOSX1
X_3253_ _3253_/A _2950_/B _3252_/Y _3201_/D gnd _3257_/B vdd OAI22X1
X_2135_ _2135_/A gnd _2137_/B vdd INVX1
X_3184_ gnd _3340_/B gnd _3184_/Y vdd NAND2X1
X_2204_ _2204_/A _2361_/A gnd _2204_/Y vdd NOR2X1
X_2899_ _2899_/A gnd _2900_/D vdd INVX1
X_2968_ _2965_/A _2965_/B gnd _2968_/Y vdd AND2X2
X_4569_ _4488_/B _4436_/CLK _4491_/Y gnd vdd DFFPOSX1
X_3871_ _3804_/A _3870_/B _3871_/C gnd _4311_/D vdd OAI21X1
X_3940_ _2406_/A _3941_/B _4162_/C gnd _3940_/Y vdd OAI21X1
X_2684_ _4017_/A _2735_/A _2110_/A _2683_/Y gnd _2684_/Y vdd OAI22X1
X_2753_ _2292_/B _2713_/A gnd _2755_/C vdd OR2X2
X_2822_ _2482_/A _2822_/B gnd _2824_/B vdd NAND2X1
X_4354_ _4354_/Q _4359_/CLK _3794_/Y gnd vdd DFFPOSX1
X_4423_ _4423_/Q _4359_/CLK _4295_/Y gnd vdd DFFPOSX1
X_4285_ _3794_/A _4283_/B _4284_/Y gnd _4285_/Y vdd AOI21X1
X_3305_ _3305_/A _2950_/B _3304_/Y _3201_/D gnd _3309_/B vdd OAI22X1
XSFILL29520x16100 gnd vdd FILL
X_3236_ gnd _3340_/B gnd _3237_/C vdd NAND2X1
X_3098_ _2471_/Y gnd _3098_/Y vdd INVX1
X_2118_ _2118_/A _4585_/B gnd _2119_/C vdd NAND2X1
X_3167_ _3167_/A _3141_/B gnd _3170_/B vdd NAND2X1
XSFILL59120x34100 gnd vdd FILL
XSFILL44080x12100 gnd vdd FILL
X_4070_ _4070_/A _4068_/Y _4004_/C _4070_/D gnd _4071_/A vdd OAI22X1
X_3021_ gnd gnd _3022_/C vdd INVX1
XSFILL59280x4100 gnd vdd FILL
X_2805_ _2456_/A _2801_/B gnd _2805_/Y vdd NOR2X1
X_3854_ _3854_/A _3852_/B gnd _3854_/Y vdd NAND2X1
X_3923_ _3922_/Y _3923_/B _3909_/C _3923_/D gnd _3928_/B vdd OAI22X1
X_2736_ _2736_/A _2736_/B _2736_/C gnd _2743_/B vdd OAI21X1
X_2667_ _2761_/A gnd _2668_/B vdd INVX1
X_4406_ _4245_/B _4417_/CLK _3695_/Y gnd vdd DFFPOSX1
X_3785_ _4153_/A _3786_/B gnd _3785_/Y vdd NAND2X1
X_4337_ _4337_/Q _4417_/CLK _3892_/Y gnd vdd DFFPOSX1
X_3219_ _3219_/A _3141_/B gnd _3222_/B vdd NAND2X1
X_4268_ _3935_/A _4269_/B gnd _4268_/Y vdd NOR2X1
X_2598_ _2418_/A gnd _2599_/D vdd INVX1
X_4199_ _4199_/A _4199_/B _4199_/C gnd _4200_/A vdd OAI21X1
XBUFX2_insert43 _4448_/Q gnd _2110_/A vdd BUFX2
XBUFX2_insert65 _2968_/Y gnd _3294_/B vdd BUFX2
XBUFX2_insert21 _3564_/Y gnd _3616_/B vdd BUFX2
XBUFX2_insert54 _4445_/Q gnd _2723_/B vdd BUFX2
XBUFX2_insert10 _3839_/Y gnd _3852_/B vdd BUFX2
XBUFX2_insert76 _4433_/Q gnd _2682_/A vdd BUFX2
XBUFX2_insert87 _3644_/Q gnd _4012_/S vdd BUFX2
XSFILL43920x42100 gnd vdd FILL
XBUFX2_insert98 _4427_/Q gnd _2895_/A vdd BUFX2
XBUFX2_insert231 _4449_/Q gnd _2922_/B vdd BUFX2
XBUFX2_insert220 _3651_/Y gnd _3683_/B vdd BUFX2
XBUFX2_insert242 _4437_/Q gnd _2330_/B vdd BUFX2
XBUFX2_insert253 _4434_/Q gnd _2676_/A vdd BUFX2
X_2521_ _2519_/Y _2520_/Y gnd _2522_/B vdd NOR2X1
XBUFX2_insert275 _4087_/Y gnd _4180_/B vdd BUFX2
XBUFX2_insert286 _4428_/Q gnd _2913_/D vdd BUFX2
XBUFX2_insert297 _4425_/Q gnd _2906_/A vdd BUFX2
X_3570_ _3570_/A _3613_/B _3570_/C gnd _3570_/Y vdd AOI21X1
XBUFX2_insert264 _4431_/Q gnd _2136_/B vdd BUFX2
XFILL71280x10100 gnd vdd FILL
X_4053_ _4231_/A _4002_/B gnd _4053_/Y vdd NOR2X1
X_2383_ _2383_/A _2383_/B _2383_/C _2382_/Y gnd _2384_/C vdd OAI22X1
X_4122_ _3944_/A _4124_/S _4111_/C gnd _4123_/A vdd OAI21X1
XSFILL29520x8100 gnd vdd FILL
X_2452_ _2609_/A _2706_/B gnd _2452_/Y vdd XNOR2X1
XSFILL14320x48100 gnd vdd FILL
X_3004_ _3004_/A _3004_/B gnd _3016_/B vdd NOR2X1
X_3837_ _3804_/A _3832_/B _3836_/Y gnd _4391_/D vdd AOI21X1
X_3768_ _3902_/A _3767_/B _3768_/C gnd _4326_/D vdd OAI21X1
X_3906_ _3773_/A _4376_/Q _3920_/S gnd _3906_/Y vdd MUX2X1
X_2719_ _2896_/A _2706_/D gnd _2719_/Y vdd NOR2X1
X_3699_ _3699_/A gnd _3771_/B vdd INVX1
XSFILL44880x8100 gnd vdd FILL
X_3622_ _3575_/A data_in[8] gnd _3624_/B vdd NAND2X1
X_2504_ _2503_/Y gnd _2504_/Y vdd INVX1
X_3484_ _3484_/A gnd _3485_/C vdd INVX1
X_2435_ _2794_/A _2434_/Y gnd _2443_/A vdd NAND2X1
X_3553_ _3553_/A gnd _3554_/B vdd INVX1
X_2366_ _2829_/B _2862_/A gnd _3271_/A vdd AND2X2
X_4036_ _4214_/A _4036_/B _4004_/C gnd _4036_/Y vdd OAI21X1
XSFILL29520x24100 gnd vdd FILL
XSFILL30000x12100 gnd vdd FILL
X_2297_ _2298_/A _2298_/B gnd _2297_/Y vdd NOR2X1
X_4105_ _4105_/A _4103_/Y _4101_/C _4102_/Y gnd _4105_/Y vdd OAI22X1
XSFILL44720x100 gnd vdd FILL
XSFILL14800x44100 gnd vdd FILL
XSFILL59120x42100 gnd vdd FILL
XSFILL44080x20100 gnd vdd FILL
XSFILL28880x52100 gnd vdd FILL
X_2082_ _2146_/Y gnd adrs_bus[10] vdd BUFX2
X_2151_ _2151_/A _4228_/A gnd _2151_/Y vdd NAND2X1
X_2220_ _2221_/B _2219_/Y gnd _3189_/A vdd XNOR2X1
X_2984_ _2984_/A _3194_/B _3194_/C gnd _2988_/A vdd NAND3X1
X_3605_ _3555_/A _3605_/B gnd _3606_/A vdd NAND2X1
X_4585_ _3562_/A _4585_/B gnd _4585_/Y vdd NAND2X1
X_3398_ _3398_/A _3396_/Y _3391_/A gnd _3401_/C vdd OAI21X1
X_3467_ _3495_/A _3466_/Y _3467_/C gnd _3467_/Y vdd NAND3X1
X_3536_ _3535_/Y _3508_/B _3508_/C gnd _3536_/Y vdd NAND3X1
X_2418_ _2418_/A _4600_/B gnd _2418_/Y vdd XNOR2X1
X_4019_ _4354_/Q _3826_/A _4074_/S gnd _4022_/D vdd MUX2X1
X_2349_ _2515_/A _2516_/A gnd _3225_/A vdd OR2X2
XSFILL43920x50100 gnd vdd FILL
X_4370_ _3726_/C _4359_/CLK _3727_/Y gnd vdd DFFPOSX1
X_3252_ gnd gnd _3252_/Y vdd INVX1
X_3321_ _3320_/Y _3321_/B gnd _3321_/Y vdd AND2X2
X_3183_ gnd gnd _3185_/A vdd INVX1
X_2203_ _2361_/B _2361_/A gnd _2213_/B vdd AND2X2
X_2134_ _2124_/A _2134_/B _2134_/C gnd _2092_/A vdd OAI21X1
X_2967_ _2967_/A _3340_/B gnd _2970_/C vdd NAND2X1
X_4568_ _4488_/A _4297_/CLK _4568_/D gnd vdd DFFPOSX1
X_2898_ _2377_/A gnd _2898_/Y vdd INVX1
X_4499_ _4501_/B gnd _4499_/Y vdd INVX1
X_3519_ _3519_/A gnd _3520_/C vdd INVX1
X_3870_ _3870_/A _3870_/B gnd _3871_/C vdd NAND2X1
X_2821_ _2817_/Y _2820_/Y _2814_/Y gnd _2825_/A vdd NAND3X1
X_2683_ _2875_/A gnd _2683_/Y vdd INVX1
X_4422_ _4292_/A _4407_/CLK _4293_/Y gnd vdd DFFPOSX1
X_2752_ _2752_/A _2711_/A gnd _2752_/Y vdd NAND2X1
X_4284_ _4418_/Q _4283_/B gnd _4284_/Y vdd NOR2X1
X_4353_ _4186_/A _4417_/CLK _4353_/D gnd vdd DFFPOSX1
X_3304_ gnd gnd _3304_/Y vdd INVX1
X_3235_ gnd gnd _3235_/Y vdd INVX1
XSFILL14480x10100 gnd vdd FILL
X_3166_ _3166_/A _3162_/Y _3165_/Y gnd _3166_/Y vdd NAND3X1
X_3097_ _3095_/Y _2950_/B _3097_/C _3201_/D gnd _3101_/B vdd OAI22X1
X_2117_ _4470_/C gnd _2119_/B vdd INVX1
X_3999_ _4320_/Q _4052_/S _4065_/C gnd _4000_/A vdd OAI21X1
XSFILL59600x28100 gnd vdd FILL
X_3020_ _2445_/Y gnd _3020_/Y vdd INVX1
X_3784_ _3717_/A _3786_/B _3784_/C gnd _3784_/Y vdd OAI21X1
X_2804_ _2104_/A _2801_/C gnd _2806_/A vdd NAND2X1
X_3853_ _3752_/A _3846_/B _3853_/C gnd _4302_/D vdd OAI21X1
X_3922_ _4313_/Q _3920_/S _3909_/C gnd _3922_/Y vdd OAI21X1
X_2735_ _2735_/A _4017_/A _2735_/C gnd _2736_/A vdd OAI21X1
X_2666_ _2665_/A _2663_/Y gnd _2670_/A vdd NAND2X1
X_4336_ _4003_/A _4373_/CLK _4336_/D gnd vdd DFFPOSX1
X_4405_ _3691_/A _4359_/CLK _4405_/D gnd vdd DFFPOSX1
X_2597_ _2312_/A gnd _2599_/A vdd INVX1
X_4198_ _3726_/C _4198_/B gnd _4198_/Y vdd NOR2X1
X_3218_ _3218_/A _3218_/B _3217_/Y gnd _3223_/A vdd NAND3X1
X_4267_ _3843_/A _4269_/B _4267_/C gnd _4267_/Y vdd AOI21X1
X_3149_ _3147_/Y _2950_/B _3149_/C _3201_/D gnd _3153_/B vdd OAI22X1
XSFILL14000x28100 gnd vdd FILL
XBUFX2_insert77 _4433_/Q gnd _4195_/A vdd BUFX2
XBUFX2_insert99 _4455_/Q gnd _2849_/A vdd BUFX2
XBUFX2_insert44 _4448_/Q gnd _2786_/C vdd BUFX2
XBUFX2_insert88 _3644_/Q gnd _4052_/S vdd BUFX2
XBUFX2_insert11 _3839_/Y gnd _3866_/B vdd BUFX2
XBUFX2_insert55 _4445_/Q gnd _2633_/B vdd BUFX2
XBUFX2_insert66 _2968_/Y gnd _3164_/B vdd BUFX2
XFILL71120x100 gnd vdd FILL
XBUFX2_insert254 _4434_/Q gnd _2516_/A vdd BUFX2
XBUFX2_insert232 _4449_/Q gnd _4017_/A vdd BUFX2
XBUFX2_insert210 _3641_/Q gnd _4241_/S vdd BUFX2
XBUFX2_insert276 _4087_/Y gnd _4231_/B vdd BUFX2
XBUFX2_insert243 _4437_/Q gnd _2574_/A vdd BUFX2
XBUFX2_insert221 _3651_/Y gnd _3685_/B vdd BUFX2
XBUFX2_insert265 _4431_/Q gnd _2915_/A vdd BUFX2
X_2520_ _2520_/A _2252_/A gnd _2520_/Y vdd AND2X2
XSFILL29040x44100 gnd vdd FILL
X_2451_ _2535_/C _2445_/B _2451_/C gnd _2451_/Y vdd AOI21X1
XBUFX2_insert287 _4428_/Q gnd _2606_/D vdd BUFX2
XBUFX2_insert298 _4425_/Q gnd _4585_/B vdd BUFX2
X_4052_ _3799_/A _4389_/Q _4052_/S gnd _4055_/D vdd MUX2X1
X_2382_ _2382_/A _2682_/A gnd _2382_/Y vdd NOR2X1
X_4121_ _4363_/Q _4158_/B gnd _4123_/B vdd NOR2X1
X_3003_ _3001_/Y _3341_/B _3003_/C gnd _3004_/B vdd OAI21X1
X_3905_ _3905_/A gnd _4027_/S vdd INVX8
X_3836_ _3836_/A _3832_/B gnd _3836_/Y vdd NOR2X1
X_3767_ _3767_/A _3767_/B gnd _3768_/C vdd NAND2X1
X_2718_ _2609_/A _2717_/B gnd _2718_/Y vdd NAND2X1
X_3698_ _3804_/A _3683_/B _3697_/Y gnd _3698_/Y vdd AOI21X1
X_2649_ _2571_/B _2571_/A gnd _2650_/B vdd NOR2X1
X_4319_ _4166_/A _4383_/CLK _3754_/Y gnd vdd DFFPOSX1
XSFILL59120x4100 gnd vdd FILL
X_3621_ _3620_/Y _3621_/B _3579_/C gnd _3633_/D vdd AOI21X1
X_3552_ _3561_/A _3552_/B gnd _3469_/B vdd NOR2X1
X_2503_ _2228_/A _2502_/B gnd _2503_/Y vdd NAND2X1
X_2365_ _2515_/A _2516_/A gnd _3245_/A vdd AND2X2
X_3483_ _3518_/A _4605_/A gnd _3483_/Y vdd NAND2X1
X_2434_ _2619_/A gnd _2434_/Y vdd INVX1
XSFILL29520x40100 gnd vdd FILL
X_4035_ _3862_/A _3932_/B gnd _4037_/B vdd NOR2X1
X_2296_ _2294_/Y _2296_/B gnd _3006_/A vdd NOR2X1
X_4104_ _4329_/Q _4098_/S _4101_/C gnd _4105_/A vdd OAI21X1
X_3819_ _3752_/A _3819_/B _3818_/Y gnd _4382_/D vdd AOI21X1
XSFILL59600x36100 gnd vdd FILL
XSFILL44560x14100 gnd vdd FILL
X_2150_ _2150_/A gnd _2152_/B vdd INVX1
X_2081_ _2081_/A gnd adrs_bus[1] vdd BUFX2
X_2983_ _2355_/Y _3141_/B gnd _2983_/Y vdd NAND2X1
XSFILL44240x2100 gnd vdd FILL
XFILL71280x16100 gnd vdd FILL
X_3604_ _3564_/A data_in[0] gnd _3606_/B vdd NAND2X1
X_3535_ data_in[15] gnd _3535_/Y vdd INVX1
XSFILL44720x8100 gnd vdd FILL
X_4584_ _4584_/A gnd _4586_/B vdd INVX1
X_2348_ _2382_/A _2682_/A gnd _3199_/A vdd OR2X2
X_3397_ _3382_/Y _3390_/B gnd _3398_/A vdd NOR2X1
X_3466_ _3465_/Y _3508_/B _3508_/C gnd _3466_/Y vdd NAND3X1
X_2417_ _2371_/A _2136_/B gnd _2417_/Y vdd XNOR2X1
X_4018_ _4018_/A _4207_/B _4017_/Y gnd _4449_/D vdd AOI21X1
X_2279_ _2232_/A _2251_/A gnd _2280_/C vdd NOR2X1
XSFILL29040x52100 gnd vdd FILL
X_3251_ _3251_/A gnd _3253_/A vdd INVX1
X_3182_ _3182_/A _3130_/B _3181_/Y _3130_/D gnd _3182_/Y vdd OAI22X1
X_3320_ gnd _3294_/B _3268_/C gnd _3320_/Y vdd NAND3X1
X_2202_ _2202_/A _2202_/B gnd _2202_/Y vdd XNOR2X1
X_2133_ _2124_/A _4600_/B gnd _2134_/C vdd NAND2X1
X_2966_ _2986_/C _2966_/B gnd _3340_/B vdd NOR2X1
X_2897_ _2895_/Y _2377_/A _2896_/Y _2406_/A gnd _2901_/A vdd AOI22X1
X_4498_ _4498_/A _4498_/B _4557_/C gnd _4498_/Y vdd AOI21X1
X_3518_ _3518_/A _4620_/A gnd _3524_/A vdd NAND2X1
X_4567_ _4476_/C _4297_/CLK _4567_/D gnd vdd DFFPOSX1
XSFILL14160x6100 gnd vdd FILL
X_3449_ _3068_/Y gnd _3449_/Y vdd INVX1
XSFILL59120x48100 gnd vdd FILL
XSFILL44080x26100 gnd vdd FILL
X_2751_ _2752_/A _2711_/A gnd _2751_/Y vdd OR2X2
X_2820_ _2820_/A _2606_/D _2823_/A gnd _2820_/Y vdd AOI21X1
X_2682_ _2682_/A gnd _2735_/A vdd INVX1
X_4421_ _4056_/A _4407_/CLK _4291_/Y gnd vdd DFFPOSX1
X_4352_ _4352_/Q _4407_/CLK _3790_/Y gnd vdd DFFPOSX1
X_4283_ _4283_/A _4283_/B _4282_/Y gnd _4283_/Y vdd AOI21X1
X_3303_ _3303_/A gnd _3305_/A vdd INVX1
X_3234_ _3234_/A _3130_/B _3233_/Y _3130_/D gnd _3238_/A vdd OAI22X1
X_3165_ _3165_/A _3163_/Y gnd _3165_/Y vdd AND2X2
X_2116_ _2118_/A _2116_/B _2116_/C gnd _2080_/A vdd OAI21X1
X_3096_ gnd gnd _3097_/C vdd INVX1
X_3998_ _4176_/A _4002_/B gnd _3998_/Y vdd NOR2X1
X_2949_ _2969_/B _2947_/A gnd _2950_/B vdd NAND2X1
X_4619_ _4621_/A _4617_/Y _4619_/C gnd _4542_/B vdd OAI21X1
XFILL70960x8100 gnd vdd FILL
XSFILL59600x44100 gnd vdd FILL
XSFILL44560x22100 gnd vdd FILL
XFILL71280x24100 gnd vdd FILL
X_3921_ _3921_/A _3921_/B gnd _3923_/B vdd NOR2X1
X_2734_ _2730_/A _2374_/A _2734_/C gnd _2736_/C vdd OAI21X1
X_3783_ _4142_/A _3786_/B gnd _3784_/C vdd NAND2X1
X_2803_ _2456_/A _2801_/B gnd _2803_/Y vdd NAND2X1
X_3852_ _4158_/A _3852_/B gnd _3853_/C vdd NAND2X1
X_2665_ _2665_/A _2663_/Y _4228_/A _2669_/B gnd _2671_/A vdd OAI22X1
X_4404_ _3688_/A _4298_/CLK _4404_/D gnd vdd DFFPOSX1
X_2596_ _2594_/Y _2482_/B _2595_/Y _2201_/B gnd _2600_/A vdd AOI22X1
X_4335_ _3992_/A _4300_/CLK _4335_/D gnd vdd DFFPOSX1
X_4197_ _4354_/Q _3826_/A _4252_/S gnd _4200_/D vdd MUX2X1
X_3217_ _3216_/Y _3215_/Y gnd _3217_/Y vdd AND2X2
X_4266_ _4266_/A _4287_/B gnd _4267_/C vdd NOR2X1
X_3148_ gnd gnd _3149_/C vdd INVX1
X_3079_ gnd gnd _3081_/A vdd INVX1
XBUFX2_insert78 _4433_/Q gnd _2874_/A vdd BUFX2
XBUFX2_insert12 _3839_/Y gnd _3870_/B vdd BUFX2
XBUFX2_insert45 _4439_/Q gnd _2283_/A vdd BUFX2
XBUFX2_insert67 _3872_/Y gnd _3893_/B vdd BUFX2
XBUFX2_insert89 _3644_/Q gnd _4030_/S vdd BUFX2
XBUFX2_insert56 _4445_/Q gnd _2307_/A vdd BUFX2
XBUFX2_insert233 _4449_/Q gnd _2382_/A vdd BUFX2
XBUFX2_insert244 _4437_/Q gnd _2772_/B vdd BUFX2
XBUFX2_insert277 _4087_/Y gnd _4198_/B vdd BUFX2
XBUFX2_insert222 _3651_/Y gnd _3680_/B vdd BUFX2
XBUFX2_insert255 _3907_/Y gnd _3932_/B vdd BUFX2
XBUFX2_insert288 _4428_/Q gnd _2127_/B vdd BUFX2
XBUFX2_insert266 _4431_/Q gnd _2346_/B vdd BUFX2
XBUFX2_insert200 _3409_/Y gnd _2118_/A vdd BUFX2
XBUFX2_insert211 _3641_/Q gnd _4153_/S vdd BUFX2
XBUFX2_insert299 _4425_/Q gnd _2295_/B vdd BUFX2
X_2381_ _4017_/A _4195_/A gnd _2383_/C vdd AND2X2
X_2450_ _2104_/A _2450_/B gnd _2451_/C vdd NOR2X1
X_4051_ _4049_/Y _4217_/B _4050_/Y gnd _4051_/Y vdd AOI21X1
X_4120_ _4347_/Q _4379_/Q _4124_/S gnd _4123_/D vdd MUX2X1
X_3002_ gnd _3340_/B gnd _3003_/C vdd NAND2X1
X_3904_ _3804_/A _3904_/B _3903_/Y gnd _3904_/Y vdd AOI21X1
XSFILL14480x16100 gnd vdd FILL
X_3697_ _4407_/Q _3683_/B gnd _3697_/Y vdd NOR2X1
X_3766_ _3692_/A _3767_/B _3765_/Y gnd _4325_/D vdd OAI21X1
XSFILL29520x38100 gnd vdd FILL
XSFILL30000x26100 gnd vdd FILL
X_2717_ _2895_/A _2717_/B gnd _2717_/Y vdd NOR2X1
X_3835_ _3902_/A _3824_/B _3835_/C gnd _3835_/Y vdd AOI21X1
X_2579_ _2673_/A _2637_/C gnd _2583_/A vdd NAND2X1
X_4249_ _4249_/A _4244_/Y _4205_/S gnd _4251_/A vdd MUX2X1
X_2648_ _2659_/A _2567_/Y gnd _2650_/A vdd NOR2X1
X_4318_ _3751_/A _4394_/CLK _4318_/D gnd vdd DFFPOSX1
XSFILL29200x20100 gnd vdd FILL
XSFILL44080x34100 gnd vdd FILL
X_2502_ _2228_/A _2502_/B gnd _2502_/Y vdd NOR2X1
X_3620_ _3553_/A _3616_/B gnd _3620_/Y vdd NAND2X1
X_3551_ _3561_/B gnd _3552_/B vdd INVX1
X_2364_ _2382_/A _2682_/A gnd _3219_/A vdd AND2X2
X_2433_ _2433_/A _2429_/A gnd _2433_/Y vdd XOR2X1
X_3482_ _3476_/Y _3481_/Y gnd _3482_/Y vdd NAND2X1
X_4103_ _4297_/Q _4158_/B gnd _4103_/Y vdd NOR2X1
X_4034_ _4212_/A _4212_/B _4036_/B gnd _4034_/Y vdd MUX2X1
X_2295_ _2295_/A _2295_/B gnd _2296_/B vdd AND2X2
X_3818_ _4153_/B _3819_/B gnd _3818_/Y vdd NOR2X1
X_3749_ _3966_/A _3754_/B gnd _3749_/Y vdd NAND2X1
XSFILL44880x48100 gnd vdd FILL
XSFILL59280x10100 gnd vdd FILL
XSFILL59600x52100 gnd vdd FILL
XSFILL44560x30100 gnd vdd FILL
X_2080_ _2080_/A gnd adrs_bus[0] vdd BUFX2
X_2982_ _2982_/A _2982_/B gnd _3141_/B vdd NOR2X1
X_3603_ _3603_/A _3603_/B _3615_/C gnd _3637_/D vdd AOI21X1
X_3465_ data_in[5] gnd _3465_/Y vdd INVX1
X_4583_ _4586_/A _4583_/B _4582_/Y gnd _4583_/Y vdd OAI21X1
X_3534_ _3513_/A _3513_/B _3534_/C gnd _3537_/C vdd OAI21X1
X_2347_ _2421_/A _4184_/A gnd _3173_/A vdd OR2X2
X_2416_ _2416_/A _2407_/Y _2416_/C gnd _2416_/Y vdd NOR3X1
X_3396_ _3384_/A _3396_/B _3396_/C _3396_/D gnd _3396_/Y vdd AOI22X1
X_2278_ _2278_/A _2278_/B _2278_/C gnd _2278_/Y vdd AOI21X1
X_4017_ _4017_/A _4207_/B _4206_/C gnd _4017_/Y vdd OAI21X1
X_3181_ gnd gnd _3181_/Y vdd INVX1
X_3250_ _3250_/A _3250_/B _3250_/C gnd _3498_/A vdd NAND3X1
X_2201_ _2204_/A _2201_/B gnd _2202_/B vdd XNOR2X1
X_2132_ _4501_/B gnd _2134_/B vdd INVX1
XSFILL29520x46100 gnd vdd FILL
XSFILL30000x34100 gnd vdd FILL
X_2965_ _2965_/A _2965_/B gnd _2986_/C vdd NAND2X1
X_2896_ _2896_/A gnd _2896_/Y vdd INVX1
XSFILL14480x24100 gnd vdd FILL
X_4497_ _4558_/B _4598_/Y _4495_/A _4556_/D gnd _4498_/B vdd AOI22X1
X_3517_ _3517_/A _3516_/Y gnd _3517_/Y vdd NAND2X1
X_4566_ _4470_/C _4297_/CLK _4566_/D gnd vdd DFFPOSX1
X_3448_ _3532_/A _3546_/Y gnd _3454_/A vdd NAND2X1
X_3379_ _3379_/A _3379_/B gnd _3380_/C vdd NOR2X1
XSFILL44080x42100 gnd vdd FILL
X_2681_ _2874_/A _2679_/Y _2681_/C _2875_/A gnd _2735_/C vdd OAI22X1
X_2750_ _2750_/A _2748_/Y gnd _2758_/C vdd NOR2X1
X_4282_ _4417_/Q _4283_/B gnd _4282_/Y vdd NOR2X1
X_4420_ _4045_/A _4298_/CLK _4289_/Y gnd vdd DFFPOSX1
X_3302_ _3302_/A _3290_/Y _3301_/Y gnd _3512_/A vdd NAND3X1
X_4351_ _4351_/Q _4345_/CLK _3788_/Y gnd vdd DFFPOSX1
X_3233_ gnd gnd _3233_/Y vdd INVX1
X_3095_ _2344_/Y gnd _3095_/Y vdd INVX1
X_2115_ _2429_/B _2118_/A gnd _2116_/C vdd NAND2X1
X_3164_ gnd _3164_/B _3164_/C gnd _3165_/A vdd NAND3X1
X_3997_ _4352_/Q _3997_/B _4052_/S gnd _3997_/Y vdd MUX2X1
X_4618_ _4621_/A _4228_/A gnd _4619_/C vdd NAND2X1
X_2948_ _2986_/B _2944_/Y gnd _2969_/B vdd NOR2X1
X_2879_ _2915_/A gnd _2879_/Y vdd INVX1
X_4549_ _4558_/B _4549_/B _4578_/Q _4556_/D gnd _4549_/Y vdd AOI22X1
XSFILL14000x6100 gnd vdd FILL
X_3851_ _3717_/A _3852_/B _3851_/C gnd _3851_/Y vdd OAI21X1
X_3920_ _4345_/Q _4377_/Q _3920_/S gnd _3923_/D vdd MUX2X1
X_2733_ _2731_/Y _2732_/Y _2733_/C gnd _2736_/B vdd NAND3X1
XFILL71280x40100 gnd vdd FILL
X_2664_ _4050_/A gnd _2669_/B vdd INVX1
X_3782_ _4273_/A _3786_/B _3781_/Y gnd _3782_/Y vdd OAI21X1
X_2802_ _2798_/Y _2801_/Y gnd _2838_/A vdd NOR2X1
X_4403_ _4212_/B _4373_/CLK _4403_/D gnd vdd DFFPOSX1
X_2595_ _2916_/A gnd _2595_/Y vdd INVX1
X_4265_ _3740_/A _4277_/B _4264_/Y gnd _4265_/Y vdd AOI21X1
X_4334_ _4334_/Q _4394_/CLK _3886_/Y gnd vdd DFFPOSX1
X_4196_ _4196_/A _4240_/B _4195_/Y gnd _4196_/Y vdd AOI21X1
X_3216_ gnd _3346_/B _3346_/C gnd _3216_/Y vdd NAND3X1
X_3147_ _2346_/Y gnd _3147_/Y vdd INVX1
X_3078_ _3076_/Y _3130_/B _3078_/C _3130_/D gnd _3082_/A vdd OAI22X1
XBUFX2_insert13 _3839_/Y gnd _3862_/B vdd BUFX2
XBUFX2_insert79 _4433_/Q gnd _2318_/B vdd BUFX2
XBUFX2_insert46 _4439_/Q gnd _2762_/A vdd BUFX2
XBUFX2_insert57 _4445_/Q gnd _2190_/B vdd BUFX2
XSFILL29200x18100 gnd vdd FILL
XBUFX2_insert68 _3872_/Y gnd _3873_/B vdd BUFX2
XBUFX2_insert201 _4451_/Q gnd _2829_/B vdd BUFX2
XBUFX2_insert212 _3641_/Q gnd _4199_/B vdd BUFX2
XBUFX2_insert245 _4437_/Q gnd _2665_/A vdd BUFX2
XBUFX2_insert223 _2975_/Y gnd _3188_/B vdd BUFX2
XBUFX2_insert256 _3907_/Y gnd _3943_/B vdd BUFX2
XBUFX2_insert278 _3645_/Q gnd _3934_/C vdd BUFX2
XBUFX2_insert267 _4431_/Q gnd _2693_/B vdd BUFX2
XBUFX2_insert289 _4428_/Q gnd _2892_/A vdd BUFX2
XBUFX2_insert234 _2972_/Y gnd _3372_/C vdd BUFX2
X_2380_ _4061_/A _4239_/A gnd _2383_/A vdd NOR2X1
X_4050_ _4050_/A _4217_/B _4228_/C gnd _4050_/Y vdd OAI21X1
X_3001_ gnd gnd _3001_/Y vdd INVX1
X_3903_ _4343_/Q _3904_/B gnd _3903_/Y vdd NOR2X1
X_3834_ _4390_/Q _3832_/B gnd _3835_/C vdd NOR2X1
X_3696_ _3538_/Y gnd _3804_/A vdd INVX4
X_2647_ _2643_/Y _2925_/B _2646_/Y gnd _2647_/Y vdd OAI21X1
X_3765_ _4232_/A _3767_/B gnd _3765_/Y vdd NAND2X1
XSFILL14480x32100 gnd vdd FILL
X_2716_ _2716_/A _2716_/B _2716_/C gnd _2716_/Y vdd AOI21X1
X_2578_ _2778_/A gnd _2637_/C vdd INVX1
X_4248_ _4248_/A _4246_/Y _4254_/C _4248_/D gnd _4249_/A vdd OAI22X1
X_4317_ _3966_/A _4383_/CLK _3750_/Y gnd vdd DFFPOSX1
X_4179_ _4416_/Q _4400_/Q _4199_/B gnd _4182_/D vdd MUX2X1
XSFILL44560x28100 gnd vdd FILL
X_2501_ _2786_/A gnd _2502_/B vdd INVX1
X_3481_ _3495_/A _3480_/Y _3481_/C gnd _3481_/Y vdd NAND3X1
X_3550_ _3562_/A _3550_/B gnd _3550_/Y vdd NOR2X1
X_4033_ _4033_/A _4033_/B _4065_/C _4030_/Y gnd _4038_/B vdd OAI22X1
X_2363_ _2421_/A _2421_/B gnd _3193_/A vdd AND2X2
X_2432_ _2416_/Y _2432_/B gnd _2952_/A vdd NAND2X1
XSFILL44240x10100 gnd vdd FILL
X_2294_ _2295_/A _2295_/B gnd _2294_/Y vdd NOR2X1
X_4102_ _4266_/A _4393_/Q _4098_/S gnd _4102_/Y vdd MUX2X1
X_3748_ _4273_/A _3754_/B _3747_/Y gnd _4316_/D vdd OAI21X1
X_3817_ _3717_/A _3819_/B _3816_/Y gnd _4381_/D vdd AOI21X1
X_3679_ _4190_/B _3680_/B gnd _3679_/Y vdd NOR2X1
X_3602_ _2965_/A _3605_/B gnd _3603_/A vdd NAND2X1
X_2981_ _2986_/A _2986_/B gnd _2982_/A vdd NAND2X1
X_2415_ _2415_/A _2415_/B _2414_/Y gnd _2416_/C vdd NAND3X1
X_3533_ _3533_/A gnd _3534_/C vdd INVX1
X_3464_ _3513_/A _3513_/B _3463_/Y gnd _3467_/C vdd OAI21X1
X_4582_ _2429_/B _4586_/A gnd _4582_/Y vdd NAND2X1
X_4016_ _4015_/Y _4011_/Y _4027_/S gnd _4018_/A vdd MUX2X1
X_3395_ _2965_/A _3382_/Y gnd _3396_/D vdd NAND2X1
X_2277_ _2277_/A _2276_/Y gnd _2278_/C vdd NAND2X1
X_2346_ _2371_/A _2346_/B gnd _2346_/Y vdd OR2X2
X_3180_ gnd gnd _3182_/A vdd INVX1
X_2200_ _2199_/Y _2188_/B _2195_/Y gnd _2202_/A vdd OAI21X1
X_2131_ _2118_/A _2131_/B _2131_/C gnd _2091_/A vdd OAI21X1
X_2964_ _2844_/Y gnd _2964_/Y vdd INVX1
X_4565_ _4565_/Q _4297_/CLK _4465_/Y gnd vdd DFFPOSX1
X_2895_ _2895_/A gnd _2895_/Y vdd INVX1
XSFILL14480x40100 gnd vdd FILL
X_4496_ _4548_/C _4495_/Y _4496_/C gnd _4498_/A vdd NAND3X1
X_3378_ _3376_/Y _3378_/B _3377_/Y gnd _3379_/B vdd NAND3X1
X_3447_ _3441_/Y _3446_/Y gnd _3447_/Y vdd NAND2X1
X_3516_ _3495_/A _3515_/Y _3516_/C gnd _3516_/Y vdd NAND3X1
X_2329_ _2329_/A _2329_/B gnd _3292_/A vdd NOR2X1
XSFILL28720x14100 gnd vdd FILL
XSFILL59280x16100 gnd vdd FILL
XSFILL44560x36100 gnd vdd FILL
X_2680_ _2110_/A gnd _2681_/C vdd INVX1
X_4281_ _4281_/A _4292_/B _4280_/Y gnd _4281_/Y vdd AOI21X1
X_3301_ _3301_/A _3300_/Y gnd _3301_/Y vdd NOR2X1
X_3232_ gnd gnd _3234_/A vdd INVX1
X_4350_ _4153_/A _4383_/CLK _3786_/Y gnd vdd DFFPOSX1
XFILL71280x38100 gnd vdd FILL
X_2114_ _4565_/Q gnd _2116_/B vdd INVX1
X_3163_ _2210_/Y _2977_/B _3090_/B gnd _3163_/Y vdd NAND3X1
X_3094_ _3075_/Y _3094_/B _3093_/Y gnd _3094_/Y vdd NAND3X1
X_2947_ _2947_/A _2946_/Y gnd _3201_/D vdd NAND2X1
X_3996_ _3996_/A _3951_/B _3995_/Y gnd _4447_/D vdd AOI21X1
X_2878_ _2878_/A _2877_/Y _2861_/Y gnd _2930_/A vdd NAND3X1
XSFILL60080x40100 gnd vdd FILL
X_4548_ _4578_/Q _4548_/B _4548_/C gnd _4548_/Y vdd OAI21X1
X_4617_ _4617_/A gnd _4617_/Y vdd INVX1
X_4479_ _4479_/A _4469_/A _4486_/A gnd _4482_/B vdd OAI21X1
XSFILL29840x4100 gnd vdd FILL
XSFILL59760x12100 gnd vdd FILL
X_3781_ _4131_/A _3786_/B gnd _3781_/Y vdd NAND2X1
X_3850_ _3969_/A _3852_/B gnd _3851_/C vdd NAND2X1
X_2801_ _2456_/A _2801_/B _2801_/C _2104_/A gnd _2801_/Y vdd OAI22X1
X_2732_ _2676_/A _2674_/D gnd _2732_/Y vdd NAND2X1
X_4402_ _3682_/A _4359_/CLK _4402_/D gnd vdd DFFPOSX1
X_2663_ _4061_/A gnd _2663_/Y vdd INVX1
X_2594_ _2915_/A gnd _2594_/Y vdd INVX1
X_4195_ _4195_/A _4240_/B _4206_/C gnd _4195_/Y vdd OAI21X1
X_3215_ _3215_/A _3345_/B _3188_/B gnd _3215_/Y vdd NAND3X1
X_4333_ _3970_/A _4300_/CLK _3884_/Y gnd vdd DFFPOSX1
X_4264_ _4408_/Q _4277_/B gnd _4264_/Y vdd NOR2X1
X_3146_ _3127_/Y _3146_/B _3145_/Y gnd _3146_/Y vdd NAND3X1
X_3077_ gnd gnd _3078_/C vdd INVX1
XBUFX2_insert14 _4450_/Q gnd _4028_/A vdd BUFX2
XBUFX2_insert47 _4439_/Q gnd _4261_/A vdd BUFX2
XBUFX2_insert36 _3738_/Y gnd _3764_/B vdd BUFX2
X_3979_ _4276_/A _4157_/B _3992_/B gnd _3982_/D vdd MUX2X1
XSFILL14160x12100 gnd vdd FILL
XBUFX2_insert58 _4445_/Q gnd _2395_/A vdd BUFX2
XBUFX2_insert69 _3872_/Y gnd _3879_/B vdd BUFX2
XBUFX2_insert202 _4451_/Q gnd _2252_/B vdd BUFX2
XBUFX2_insert213 _3641_/Q gnd _4245_/S vdd BUFX2
XBUFX2_insert224 _2975_/Y gnd _3194_/B vdd BUFX2
XBUFX2_insert257 _3907_/Y gnd _4002_/B vdd BUFX2
XBUFX2_insert246 _4437_/Q gnd _4239_/A vdd BUFX2
XBUFX2_insert268 _4431_/Q gnd _2482_/A vdd BUFX2
XBUFX2_insert279 _3645_/Q gnd _3988_/C vdd BUFX2
XBUFX2_insert235 _2972_/Y gnd _3164_/C vdd BUFX2
X_3000_ _2998_/Y _3130_/B _3000_/C _3130_/D gnd _3004_/A vdd OAI22X1
X_3902_ _3902_/A _3893_/B _3901_/Y gnd _4342_/D vdd AOI21X1
X_3764_ _3764_/A _3764_/B _3763_/Y gnd _3764_/Y vdd OAI21X1
X_3833_ _3692_/A _3832_/B _3832_/Y gnd _3833_/Y vdd AOI21X1
X_2577_ _2577_/A _2577_/B gnd _2577_/Y vdd NOR2X1
X_2646_ _2574_/A _2646_/B _2745_/A _2645_/Y gnd _2646_/Y vdd OAI22X1
X_3695_ _3902_/A _3680_/B _3694_/Y gnd _3695_/Y vdd AOI21X1
XSFILL14960x2100 gnd vdd FILL
X_2715_ _2392_/B _2715_/B gnd _2716_/B vdd NAND2X1
X_4247_ _4069_/A _4245_/S _4247_/C gnd _4248_/A vdd OAI21X1
X_4178_ _4178_/A _4176_/Y _4243_/C _4175_/Y gnd _4178_/Y vdd OAI22X1
X_4316_ _4133_/A _4300_/CLK _4316_/D gnd vdd DFFPOSX1
X_3129_ gnd gnd _3129_/Y vdd INVX1
XSFILL59280x24100 gnd vdd FILL
XFILL71280x4100 gnd vdd FILL
XSFILL44560x44100 gnd vdd FILL
X_2500_ _2500_/A _2500_/B _2496_/Y gnd _2500_/Y vdd OAI21X1
X_2431_ _2419_/Y _2431_/B _2431_/C gnd _2432_/B vdd NOR3X1
X_3480_ _3480_/A _3508_/B _3508_/C gnd _3480_/Y vdd NAND3X1
XFILL71280x46100 gnd vdd FILL
X_4032_ _4032_/A _4052_/S _4065_/C gnd _4033_/A vdd OAI21X1
X_2293_ _2293_/A _2292_/Y gnd _2293_/Y vdd NOR2X1
X_2362_ _2371_/A _2136_/B gnd _3167_/A vdd AND2X2
X_4101_ _4101_/A _4101_/B _4101_/C _4101_/D gnd _4106_/B vdd OAI22X1
X_3747_ _4133_/A _3754_/B gnd _3747_/Y vdd NAND2X1
X_3816_ _3816_/A _3819_/B gnd _3816_/Y vdd NOR2X1
X_3678_ _3496_/Y gnd _4283_/A vdd INVX4
X_2629_ _2629_/A _2627_/Y _2629_/C gnd _2629_/Y vdd OAI21X1
XSFILL44880x100 gnd vdd FILL
XSFILL59760x20100 gnd vdd FILL
X_2980_ _2980_/A _2976_/Y _2980_/C gnd _2980_/Y vdd NAND3X1
X_3601_ _3601_/A data_in[15] gnd _3603_/B vdd NAND2X1
X_4581_ _3422_/A gnd _4583_/B vdd INVX1
X_3394_ _2965_/B _3393_/Y gnd _3396_/C vdd NOR2X1
X_2414_ _2411_/Y _2410_/Y _2414_/C _2414_/D gnd _2414_/Y vdd AOI22X1
X_3463_ _3463_/A gnd _3463_/Y vdd INVX1
X_3532_ _3532_/A _4626_/A gnd _3538_/A vdd NAND2X1
X_4015_ _4014_/Y _4015_/B _4010_/C _4015_/D gnd _4015_/Y vdd OAI22X1
XSFILL14480x38100 gnd vdd FILL
X_2276_ _2202_/B _2276_/B gnd _2276_/Y vdd NOR2X1
X_2345_ _2361_/A _2361_/B gnd _3121_/A vdd OR2X2
X_2130_ _2118_/A _4597_/B gnd _2131_/C vdd NAND2X1
X_2963_ _2963_/A _3130_/B _2959_/Y _3130_/D gnd _2971_/A vdd OAI22X1
XSFILL44240x16100 gnd vdd FILL
X_4564_ _4563_/Y _4558_/Y _4557_/C gnd _4564_/Y vdd AOI21X1
X_2894_ _2919_/B _2894_/B gnd _2920_/B vdd NOR2X1
X_3515_ _3515_/A _3508_/B _3508_/C gnd _3515_/Y vdd NAND3X1
X_2328_ _2856_/A _2745_/A gnd _2329_/B vdd AND2X2
X_4495_ _4495_/A _4495_/B gnd _4495_/Y vdd NAND2X1
X_3377_ _3143_/A gnd gnd _3143_/D gnd _3377_/Y vdd AOI22X1
X_3446_ _3495_/A _3445_/Y _3443_/Y gnd _3446_/Y vdd NAND3X1
X_2259_ _2255_/Y _2259_/B gnd _3293_/A vdd XOR2X1
XSFILL59280x32100 gnd vdd FILL
XSFILL44560x52100 gnd vdd FILL
X_4280_ _4416_/Q _4292_/B gnd _4280_/Y vdd NOR2X1
X_3300_ _3298_/Y _3300_/B _3299_/Y gnd _3300_/Y vdd NAND3X1
X_3231_ _3231_/A _3231_/B gnd _3250_/A vdd NOR2X1
X_3162_ _2314_/Y _3090_/B _3110_/C gnd _3162_/Y vdd NAND3X1
X_2113_ _2113_/A gnd mem_wr vdd BUFX2
X_3093_ _3088_/Y _3093_/B gnd _3093_/Y vdd NOR2X1
X_2877_ _2922_/C _2876_/Y gnd _2877_/Y vdd NOR2X1
X_2946_ _2966_/B gnd _2946_/Y vdd INVX1
X_3995_ _2371_/A _3951_/B _3951_/C gnd _3995_/Y vdd OAI21X1
X_4547_ _4545_/Y _4547_/B gnd _4547_/Y vdd NOR2X1
X_4616_ _4612_/A _4614_/Y _4616_/C gnd _4616_/Y vdd OAI21X1
X_4478_ _4488_/A gnd _4486_/A vdd INVX2
XSFILL59440x100 gnd vdd FILL
X_3429_ _2986_/A _2986_/B gnd _3508_/B vdd NOR2X1
X_2731_ _2374_/B _2731_/B gnd _2731_/Y vdd NAND2X1
X_2800_ _2614_/C gnd _2801_/C vdd INVX1
X_3780_ _3813_/A _3802_/B _3780_/C gnd _3780_/Y vdd OAI21X1
X_4401_ _4190_/B _4417_/CLK _4401_/D gnd vdd DFFPOSX1
X_2662_ _2657_/Y _2659_/Y _2662_/C gnd _2662_/Y vdd NAND3X1
X_2593_ _2592_/Y gnd _2593_/Y vdd INVX1
X_4332_ _3881_/A _4394_/CLK _4332_/D gnd vdd DFFPOSX1
X_4194_ _4194_/A _4189_/Y _4205_/S gnd _4196_/A vdd MUX2X1
X_3214_ _3214_/A _3188_/B _3188_/C gnd _3218_/B vdd NAND3X1
X_3145_ _3140_/Y _3145_/B gnd _3145_/Y vdd NOR2X1
X_4263_ _3703_/Y _3651_/B gnd _4263_/Y vdd AND2X2
XSFILL14480x46100 gnd vdd FILL
X_3076_ gnd gnd _3076_/Y vdd INVX1
XBUFX2_insert15 _4450_/Q gnd _2098_/A vdd BUFX2
X_2929_ _2861_/Y _2929_/B _2929_/C gnd _2930_/C vdd AOI21X1
XBUFX2_insert59 _4436_/Q gnd _2745_/A vdd BUFX2
XBUFX2_insert48 _4439_/Q gnd _2659_/A vdd BUFX2
X_3978_ _3978_/A _3978_/B _3909_/C _3975_/Y gnd _3983_/B vdd OAI22X1
XBUFX2_insert37 _3738_/Y gnd _3740_/B vdd BUFX2
XBUFX2_insert203 _4451_/Q gnd _2374_/A vdd BUFX2
XBUFX2_insert236 _2972_/Y gnd _3346_/C vdd BUFX2
XBUFX2_insert258 _3907_/Y gnd _3921_/B vdd BUFX2
XBUFX2_insert247 _4443_/Q gnd _2456_/A vdd BUFX2
XBUFX2_insert225 _2975_/Y gnd _3032_/B vdd BUFX2
XBUFX2_insert214 _2943_/Y gnd _3110_/C vdd BUFX2
XBUFX2_insert269 _2960_/Y gnd _2977_/B vdd BUFX2
X_3901_ _4069_/A _3893_/B gnd _3901_/Y vdd NOR2X1
XFILL71280x100 gnd vdd FILL
X_3694_ _4245_/B _3680_/B gnd _3694_/Y vdd NOR2X1
X_3763_ _4221_/A _3764_/B gnd _3763_/Y vdd NAND2X1
X_3832_ _4389_/Q _3832_/B gnd _3832_/Y vdd NOR2X1
X_2714_ _2292_/B _2714_/B gnd _2716_/A vdd NAND2X1
X_2576_ _2574_/Y _2576_/B gnd _2577_/A vdd NAND2X1
X_2645_ _2856_/A gnd _2645_/Y vdd INVX1
X_4315_ _3944_/A _4394_/CLK _4315_/D gnd vdd DFFPOSX1
X_4246_ _4246_/A _4180_/B gnd _4246_/Y vdd NOR2X1
X_4177_ _4320_/Q _4241_/S _4243_/C gnd _4178_/A vdd OAI21X1
XSFILL29680x22100 gnd vdd FILL
X_3128_ gnd gnd _3130_/A vdd INVX1
XSFILL60080x46100 gnd vdd FILL
X_3059_ _2177_/Y _3007_/B _3032_/B gnd _3059_/Y vdd NAND3X1
XSFILL14960x42100 gnd vdd FILL
XSFILL29360x4100 gnd vdd FILL
XSFILL59760x18100 gnd vdd FILL
X_2430_ _2428_/Y _2429_/Y _2430_/C gnd _2431_/C vdd NAND3X1
X_2361_ _2361_/A _2361_/B gnd _2361_/Y vdd AND2X2
X_4031_ _4031_/A _3932_/B gnd _4033_/B vdd NOR2X1
X_2292_ _2290_/B _2292_/B gnd _2292_/Y vdd AND2X2
XSFILL43760x12100 gnd vdd FILL
X_4100_ _4313_/Q _4098_/S _4111_/C gnd _4101_/A vdd OAI21X1
X_3677_ _4281_/A _3680_/B _3676_/Y gnd _3677_/Y vdd AOI21X1
X_3746_ _3813_/A _3740_/B _3746_/C gnd _4315_/D vdd OAI21X1
X_3815_ _4273_/A _3819_/B _3815_/C gnd _4380_/D vdd AOI21X1
X_4229_ _4227_/Y _4217_/B _4228_/Y gnd _4229_/Y vdd AOI21X1
X_2559_ _2551_/Y _2558_/Y _2553_/Y gnd _2559_/Y vdd OAI21X1
XSFILL30000x2100 gnd vdd FILL
X_2628_ _2609_/A _2612_/Y gnd _2629_/C vdd NAND2X1
XSFILL14160x18100 gnd vdd FILL
XSFILL14800x2100 gnd vdd FILL
X_4580_ _2159_/A _4436_/CLK _4564_/Y gnd vdd DFFPOSX1
X_3531_ _3531_/A _3530_/Y gnd _3531_/Y vdd NAND2X1
X_3600_ _3600_/A _3598_/Y _3615_/C gnd _3636_/D vdd AOI21X1
X_3393_ _2986_/A gnd _3393_/Y vdd INVX1
X_2344_ _2395_/A _2394_/B gnd _2344_/Y vdd OR2X2
X_2413_ _2932_/B _4585_/B gnd _2414_/D vdd OR2X2
X_3462_ _3434_/A _3550_/Y gnd _3468_/A vdd NAND2X1
X_4014_ _4337_/Q _4012_/S _4010_/C gnd _4014_/Y vdd OAI21X1
XFILL71120x4100 gnd vdd FILL
X_2275_ _2346_/B _2312_/A gnd _2276_/B vdd XNOR2X1
XSFILL14960x8100 gnd vdd FILL
X_3729_ _3729_/A _3737_/B _3728_/Y gnd _4371_/D vdd OAI21X1
XSFILL14640x14100 gnd vdd FILL
X_2962_ _2961_/A _2969_/B gnd _3130_/B vdd NAND2X1
X_2893_ _2890_/Y _2892_/Y _2893_/C gnd _2894_/B vdd NAND3X1
XSFILL44240x32100 gnd vdd FILL
X_4563_ _4462_/A _4560_/Y _4562_/Y gnd _4563_/Y vdd NAND3X1
X_4494_ _4486_/A _4485_/Y _4486_/B gnd _4495_/B vdd NOR3X1
X_3514_ data_in[12] gnd _3515_/A vdd INVX1
X_3445_ _3444_/Y _3508_/B _3508_/C gnd _3445_/Y vdd NAND3X1
X_2327_ _2856_/A _2745_/A gnd _2329_/A vdd NOR2X1
X_2258_ _2257_/Y _2256_/Y gnd _2259_/B vdd NOR2X1
X_3376_ gnd _3240_/B _3324_/C gnd _3376_/Y vdd NAND3X1
XSFILL29680x30100 gnd vdd FILL
X_2189_ _2190_/A _2395_/A gnd _2191_/A vdd NAND2X1
XSFILL59760x26100 gnd vdd FILL
X_3230_ _3230_/A _3204_/B _3229_/Y _3204_/D gnd _3231_/A vdd OAI22X1
X_2112_ _2112_/A gnd mem_rd vdd BUFX2
X_3161_ gnd _3343_/B gnd _3166_/A vdd NAND2X1
X_3092_ _3090_/Y _3092_/B _3092_/C gnd _3093_/B vdd NAND3X1
X_2876_ _2922_/A _2922_/B _2876_/C gnd _2876_/Y vdd OAI21X1
X_4615_ _4612_/A _4217_/A gnd _4616_/C vdd NAND2X1
X_2945_ _2986_/B _2944_/Y gnd _2966_/B vdd NAND2X1
X_3994_ _3993_/Y _3994_/B _4027_/S gnd _3996_/A vdd MUX2X1
X_4546_ _2147_/A _2150_/A _4534_/Y gnd _4547_/B vdd NAND3X1
X_4477_ _4477_/A _4477_/B _4557_/C gnd _4567_/D vdd AOI21X1
X_3428_ data_in[0] gnd _3428_/Y vdd INVX1
X_3359_ gnd gnd _3359_/Y vdd INVX1
XSFILL14160x26100 gnd vdd FILL
X_2730_ _2730_/A _2374_/A _2677_/C _4028_/A gnd _2733_/C vdd AOI22X1
X_2661_ _2661_/A _2660_/Y gnd _2662_/C vdd NAND2X1
X_4400_ _4400_/Q _4359_/CLK _3677_/Y gnd vdd DFFPOSX1
X_4262_ _4262_/A _4240_/B _4261_/Y gnd _4439_/D vdd AOI21X1
X_2592_ _2577_/Y _2592_/B gnd _2592_/Y vdd NAND2X1
X_4331_ _3948_/A _4298_/CLK _4331_/D gnd vdd DFFPOSX1
X_4193_ _4192_/Y _4193_/B _4254_/C _4193_/D gnd _4194_/A vdd OAI22X1
X_3213_ gnd _3343_/B gnd _3218_/A vdd NAND2X1
X_3075_ _3074_/Y _3071_/Y gnd _3075_/Y vdd NOR2X1
X_3144_ _3144_/A _3141_/Y _3143_/Y gnd _3145_/B vdd NAND3X1
X_3977_ _3751_/A _3920_/S _3909_/C gnd _3978_/A vdd OAI21X1
XBUFX2_insert16 _4450_/Q gnd _2673_/A vdd BUFX2
XBUFX2_insert38 _3738_/Y gnd _3760_/B vdd BUFX2
X_2928_ _2852_/Y _2925_/Y _2927_/Y gnd _2929_/C vdd OAI21X1
X_2859_ _2772_/B _2859_/B gnd _2859_/Y vdd NAND2X1
XBUFX2_insert49 _3805_/Y gnd _3824_/B vdd BUFX2
X_4529_ _4548_/C _4540_/C _4529_/C gnd _4529_/Y vdd NAND3X1
XBUFX2_insert204 _4451_/Q gnd _4039_/A vdd BUFX2
XBUFX2_insert259 _3907_/Y gnd _4020_/B vdd BUFX2
XSFILL59280x38100 gnd vdd FILL
XBUFX2_insert237 _2972_/Y gnd _3268_/C vdd BUFX2
XBUFX2_insert226 _2975_/Y gnd _3240_/B vdd BUFX2
XBUFX2_insert248 _4443_/Q gnd _2706_/B vdd BUFX2
XBUFX2_insert215 _2943_/Y gnd _2947_/A vdd BUFX2
XSFILL14640x22100 gnd vdd FILL
X_3900_ _3692_/A _3904_/B _3899_/Y gnd _3900_/Y vdd AOI21X1
X_3831_ _3764_/A _3824_/B _3830_/Y gnd _4388_/D vdd AOI21X1
X_2644_ _2925_/B gnd _2646_/B vdd INVX1
XSFILL44240x40100 gnd vdd FILL
X_3762_ _3729_/A _3764_/B _3761_/Y gnd _4323_/D vdd OAI21X1
X_3693_ _3531_/Y gnd _3902_/A vdd INVX4
X_2713_ _2713_/A gnd _2714_/B vdd INVX1
X_2575_ _2768_/A _2100_/A gnd _2576_/B vdd XNOR2X1
X_4245_ _4292_/A _4245_/B _4245_/S gnd _4248_/D vdd MUX2X1
X_4314_ _4314_/Q _4373_/CLK _3744_/Y gnd vdd DFFPOSX1
X_4176_ _4176_/A _4231_/B gnd _4176_/Y vdd NOR2X1
X_3127_ _3126_/Y _3127_/B gnd _3127_/Y vdd NOR2X1
X_3058_ _2302_/Y _3032_/B _2947_/A gnd _3062_/B vdd NAND3X1
XSFILL44720x18100 gnd vdd FILL
X_2291_ _2290_/B _2433_/A gnd _2293_/A vdd NOR2X1
X_2360_ _2307_/A _4597_/B gnd _2360_/Y vdd AND2X2
XSFILL60240x22100 gnd vdd FILL
X_4030_ _4208_/A _4208_/B _4030_/S gnd _4030_/Y vdd MUX2X1
X_3814_ _3814_/A _3819_/B gnd _3815_/C vdd NOR2X1
X_3676_ _4400_/Q _3680_/B gnd _3676_/Y vdd NOR2X1
X_3745_ _3944_/A _3764_/B gnd _3746_/C vdd NAND2X1
X_2627_ _2614_/C _2613_/Y gnd _2627_/Y vdd NOR2X1
X_4228_ _4228_/A _4217_/B _4228_/C gnd _4228_/Y vdd OAI21X1
X_2558_ _2558_/A _2528_/Y _2557_/Y gnd _2558_/Y vdd AOI21X1
X_2489_ _2482_/A gnd _2490_/B vdd INVX1
X_4159_ _4334_/Q _4098_/S _4101_/C gnd _4159_/Y vdd OAI21X1
X_3461_ _3455_/Y _3461_/B gnd _3461_/Y vdd NAND2X1
X_3530_ _3495_/A _3529_/Y _3527_/Y gnd _3530_/Y vdd NAND3X1
X_4013_ _4191_/A _4020_/B gnd _4015_/B vdd NOR2X1
X_3392_ _2965_/A gnd _3396_/B vdd INVX1
X_2274_ _2185_/B _2191_/Y gnd _2277_/A vdd NOR2X1
X_2343_ _2428_/A _2892_/A gnd _2343_/Y vdd OR2X2
X_2412_ _2932_/B _4585_/B gnd _2414_/C vdd NAND2X1
XSFILL29680x28100 gnd vdd FILL
XSFILL45200x38100 gnd vdd FILL
X_3728_ _3732_/A _3726_/B _4031_/A gnd _3728_/Y vdd OAI21X1
X_3659_ _3811_/A _3658_/B _3659_/C gnd _3659_/Y vdd AOI21X1
XSFILL29360x10100 gnd vdd FILL
XSFILL14640x30100 gnd vdd FILL
XSFILL44560x4100 gnd vdd FILL
X_2961_ _2961_/A _2946_/Y gnd _3130_/D vdd NAND2X1
X_2892_ _2892_/A _2913_/C gnd _2892_/Y vdd NAND2X1
X_4562_ _4462_/B _2159_/A _4562_/C gnd _4562_/Y vdd NAND3X1
X_4493_ _4485_/Y _4493_/B _4493_/C gnd _4496_/C vdd OAI21X1
X_3513_ _3513_/A _3513_/B _3513_/C gnd _3516_/C vdd OAI21X1
X_3444_ data_in[2] gnd _3444_/Y vdd INVX1
X_2257_ _2351_/B _2351_/A gnd _2257_/Y vdd NOR2X1
X_2326_ _2324_/Y _2326_/B gnd _3266_/A vdd NOR2X1
X_3375_ _3375_/A _3141_/B gnd _3378_/B vdd NAND2X1
X_2188_ _2196_/A _2188_/B _2188_/C gnd _2192_/A vdd OAI21X1
XSFILL60240x30100 gnd vdd FILL
XSFILL14800x8100 gnd vdd FILL
X_2111_ _4017_/A gnd data_out[9] vdd BUFX2
X_3160_ _3160_/A _3160_/B gnd _3172_/B vdd NOR2X1
X_3091_ _3143_/A gnd gnd _3143_/D gnd _3092_/C vdd AOI22X1
X_3993_ _3992_/Y _3993_/B _3982_/C _3993_/D gnd _3993_/Y vdd OAI22X1
X_2875_ _2875_/A _2875_/B gnd _2876_/C vdd NAND2X1
X_4545_ _4578_/Q gnd _4545_/Y vdd INVX1
X_2944_ _2986_/A gnd _2944_/Y vdd INVX1
XSFILL14480x8100 gnd vdd FILL
X_4614_ _4614_/A gnd _4614_/Y vdd INVX1
X_3358_ _3358_/A gnd _3360_/A vdd INVX1
X_4476_ _4558_/B _4589_/Y _4476_/C _4556_/D gnd _4477_/A vdd AOI22X1
X_3427_ _3513_/A _3513_/B _3427_/C gnd _3427_/Y vdd OAI21X1
X_3289_ _3287_/Y _3341_/B _3289_/C gnd _3289_/Y vdd OAI21X1
X_2309_ _2361_/A _2361_/B gnd _2311_/A vdd NOR2X1
XFILL70960x16100 gnd vdd FILL
X_2660_ _2762_/C gnd _2660_/Y vdd INVX2
X_2591_ _2591_/A _2591_/B gnd _2592_/B vdd NOR2X1
X_4261_ _4261_/A _4240_/B _4239_/C gnd _4261_/Y vdd OAI21X1
X_3212_ _3212_/A _3211_/Y gnd _3212_/Y vdd NOR2X1
X_4330_ _3877_/A _4373_/CLK _4330_/D gnd vdd DFFPOSX1
X_4192_ _4337_/Q _4199_/B _4254_/C gnd _4192_/Y vdd OAI21X1
X_3074_ _3072_/Y _3204_/B _3074_/C _3204_/D gnd _3074_/Y vdd OAI22X1
X_3143_ _3143_/A gnd gnd _3143_/D gnd _3143_/Y vdd AOI22X1
X_2927_ _2848_/B _2848_/A _2927_/C gnd _2927_/Y vdd AOI21X1
X_3976_ _4366_/Q _3921_/B gnd _3978_/B vdd NOR2X1
XBUFX2_insert17 _4450_/Q gnd _2515_/A vdd BUFX2
X_2789_ _2789_/A _2788_/Y gnd _2789_/Y vdd NOR2X1
X_2858_ _2925_/B gnd _2859_/B vdd INVX1
X_4528_ _4528_/A _4528_/B _4534_/B gnd _4529_/C vdd OAI21X1
XSFILL29680x36100 gnd vdd FILL
XBUFX2_insert39 _3738_/Y gnd _3754_/B vdd BUFX2
X_4459_ _4560_/A _4458_/Y gnd _4548_/C vdd NOR2X1
XSFILL28720x52100 gnd vdd FILL
XBUFX2_insert205 _4451_/Q gnd _2779_/B vdd BUFX2
XBUFX2_insert216 _2943_/Y gnd _3188_/C vdd BUFX2
XBUFX2_insert227 _2975_/Y gnd _3267_/C vdd BUFX2
XBUFX2_insert249 _4443_/Q gnd _2301_/A vdd BUFX2
XBUFX2_insert238 _4446_/Q gnd _2361_/A vdd BUFX2
X_3761_ _4032_/A _3764_/B gnd _3761_/Y vdd NAND2X1
X_3830_ _4041_/B _3824_/B gnd _3830_/Y vdd NOR2X1
X_3692_ _3692_/A _3683_/B _3691_/Y gnd _4405_/D vdd AOI21X1
X_2574_ _2574_/A _2925_/B gnd _2574_/Y vdd XNOR2X1
X_2643_ _2574_/A gnd _2643_/Y vdd INVX1
X_2712_ _2392_/B _2715_/B gnd _2716_/C vdd NOR2X1
X_4244_ _4244_/A _4242_/Y _4243_/C _4244_/D gnd _4244_/Y vdd OAI22X1
X_4175_ _4352_/Q _3997_/B _4241_/S gnd _4175_/Y vdd MUX2X1
X_4313_ _4313_/Q _4345_/CLK _3742_/Y gnd vdd DFFPOSX1
XSFILL59440x14100 gnd vdd FILL
X_3126_ _3124_/Y _3204_/B _3125_/Y _3204_/D gnd _3126_/Y vdd OAI22X1
X_3057_ gnd _3343_/B gnd _3057_/Y vdd NAND2X1
X_3959_ _3881_/A _3968_/S _3982_/C gnd _3960_/A vdd OAI21X1
XSFILL59760x50100 gnd vdd FILL
X_2290_ _2433_/A _2290_/B gnd _2290_/Y vdd XOR2X1
X_3744_ _3811_/A _3764_/B _3743_/Y gnd _3744_/Y vdd OAI21X1
X_3813_ _3813_/A _3824_/B _3812_/Y gnd _3813_/Y vdd AOI21X1
X_2557_ _2552_/B gnd _2557_/Y vdd INVX1
X_3675_ _3489_/Y gnd _4281_/A vdd INVX4
X_2626_ _2799_/A _2612_/Y gnd _2629_/A vdd NOR2X1
X_4227_ _4226_/Y _4227_/B _4205_/S gnd _4227_/Y vdd MUX2X1
X_2488_ _2488_/A _2488_/B _2488_/C gnd _2492_/B vdd OAI21X1
X_4158_ _4158_/A _4158_/B gnd _4158_/Y vdd NOR2X1
X_4089_ _4312_/Q _4153_/S _4155_/C gnd _4090_/A vdd OAI21X1
X_3109_ gnd _3343_/B gnd _3114_/A vdd NAND2X1
XSFILL14160x50100 gnd vdd FILL
X_3391_ _3391_/A _3390_/Y gnd _3401_/A vdd NAND2X1
X_2411_ _2307_/A _2190_/A gnd _2411_/Y vdd OR2X2
X_3460_ _3495_/A _3459_/Y _3460_/C gnd _3461_/B vdd NAND3X1
X_4012_ _4417_/Q _4190_/B _4012_/S gnd _4015_/D vdd MUX2X1
X_2273_ _2287_/B _2272_/Y gnd _3345_/A vdd XNOR2X1
XSFILL29200x100 gnd vdd FILL
XSFILL14320x10100 gnd vdd FILL
X_2342_ _2301_/A _2301_/B gnd _2342_/Y vdd OR2X2
XSFILL44240x46100 gnd vdd FILL
X_3727_ _3794_/A _3737_/B _3726_/Y gnd _3727_/Y vdd OAI21X1
X_3658_ _3935_/B _3658_/B gnd _3659_/C vdd NOR2X1
X_3589_ _3589_/A data_in[11] gnd _3589_/Y vdd NAND2X1
X_2609_ _2609_/A gnd _2609_/Y vdd INVX1
X_2960_ _2965_/A _2965_/B gnd _2960_/Y vdd NOR2X1
X_4561_ _4545_/Y _4553_/Y _4547_/B gnd _4562_/C vdd NOR3X1
X_2891_ _2891_/A gnd _2913_/C vdd INVX1
X_3374_ _3369_/Y _3374_/B _3374_/C gnd _3379_/A vdd NAND3X1
X_4492_ _4495_/A gnd _4493_/C vdd INVX1
X_3512_ _3512_/A gnd _3513_/C vdd INVX1
X_3443_ _3513_/A _3513_/B _3442_/Y gnd _3443_/Y vdd OAI21X1
X_2256_ _2745_/A _2856_/A gnd _2256_/Y vdd AND2X2
X_2325_ _4039_/A _4217_/A gnd _2326_/B vdd AND2X2
X_2187_ _2187_/A _2193_/B gnd _2196_/A vdd NOR2X1
X_2110_ _2110_/A gnd data_out[8] vdd BUFX2
X_3090_ gnd _3090_/B _3116_/C gnd _3090_/Y vdd NAND3X1
X_2943_ _2982_/B gnd _2943_/Y vdd INVX8
X_3992_ _3992_/A _3992_/B _3982_/C gnd _3992_/Y vdd OAI21X1
X_2874_ _2874_/A gnd _2922_/A vdd INVX1
X_4544_ _4543_/Y _4228_/C gnd _4544_/Y vdd AND2X2
X_4613_ _4612_/A _4611_/Y _4613_/C gnd _4530_/B vdd OAI21X1
XSFILL58960x10100 gnd vdd FILL
X_3357_ _3357_/A _2950_/B _3356_/Y _3201_/D gnd _3361_/B vdd OAI22X1
X_4475_ _4548_/C _4486_/B _4475_/C gnd _4477_/B vdd NAND3X1
X_2308_ _2306_/Y _2307_/Y gnd _2308_/Y vdd NOR2X1
X_3426_ _2965_/A _2965_/B gnd _3513_/A vdd NAND2X1
X_2239_ _2252_/A gnd _2253_/A vdd INVX1
X_3288_ gnd _3340_/B gnd _3289_/C vdd NAND2X1
XSFILL44400x4100 gnd vdd FILL
XSFILL14640x36100 gnd vdd FILL
XSFILL44080x4100 gnd vdd FILL
X_2590_ _2590_/A _2642_/C _2590_/C gnd _2591_/A vdd NAND3X1
X_4191_ _4191_/A _4198_/B gnd _4193_/B vdd NOR2X1
X_4260_ _4260_/A _4260_/B _4205_/S gnd _4262_/A vdd MUX2X1
X_3211_ _3211_/A _3341_/B _3210_/Y gnd _3211_/Y vdd OAI21X1
X_3142_ gnd _3090_/B _3116_/C gnd _3144_/A vdd NAND3X1
X_3073_ gnd gnd _3074_/C vdd INVX1
X_2926_ _2762_/A _2926_/B _2846_/Y gnd _2927_/C vdd AOI21X1
X_2857_ _2768_/A _2924_/C gnd _2857_/Y vdd NAND2X1
XBUFX2_insert18 _3564_/Y gnd _3590_/B vdd BUFX2
X_3975_ _4153_/A _4153_/B _3920_/S gnd _3975_/Y vdd MUX2X1
X_2788_ _2788_/A _2787_/Y gnd _2788_/Y vdd NAND2X1
X_4527_ _4575_/Q gnd _4534_/B vdd INVX1
X_4458_ _4462_/A gnd _4458_/Y vdd INVX1
X_4389_ _4389_/Q _4407_/CLK _3833_/Y gnd vdd DFFPOSX1
X_3409_ _3387_/B _3389_/Y _3410_/B gnd _3409_/Y vdd AOI21X1
XBUFX2_insert206 _3641_/Q gnd _4098_/S vdd BUFX2
XBUFX2_insert217 _2943_/Y gnd _3292_/C vdd BUFX2
XBUFX2_insert239 _4446_/Q gnd _2201_/B vdd BUFX2
XSFILL44400x14100 gnd vdd FILL
XBUFX2_insert228 _2975_/Y gnd _3090_/B vdd BUFX2
XSFILL29840x12100 gnd vdd FILL
XFILL71120x16100 gnd vdd FILL
X_3760_ _3794_/A _3760_/B _3759_/Y gnd _4322_/D vdd OAI21X1
X_2711_ _2711_/A gnd _2715_/B vdd INVX1
X_2642_ _2637_/Y _2642_/B _2642_/C _2641_/Y gnd _2652_/B vdd OAI22X1
X_3691_ _3691_/A _3683_/B gnd _3691_/Y vdd NOR2X1
X_2573_ _2573_/A _2573_/B _2573_/C gnd _2577_/B vdd NAND3X1
X_4312_ _4312_/Q _4345_/CLK _4312_/D gnd vdd DFFPOSX1
XSFILL43760x42100 gnd vdd FILL
X_4243_ _3767_/A _4241_/S _4243_/C gnd _4244_/A vdd OAI21X1
X_4174_ _4174_/A _3951_/B _4173_/Y gnd _4431_/D vdd AOI21X1
X_3125_ gnd gnd _3125_/Y vdd INVX1
X_3056_ _3056_/A _3056_/B gnd _3068_/B vdd NOR2X1
X_3889_ _4003_/A _3896_/B gnd _3889_/Y vdd NOR2X1
X_2909_ _2896_/A _2900_/D gnd _2909_/Y vdd NOR2X1
X_3958_ _4300_/Q _3943_/B gnd _3960_/B vdd NOR2X1
X_3743_ _4314_/Q _3764_/B gnd _3743_/Y vdd NAND2X1
X_3812_ _4379_/Q _3824_/B gnd _3812_/Y vdd NOR2X1
X_3674_ _3788_/A _3671_/B _3673_/Y gnd _4399_/D vdd AOI21X1
X_2556_ _2572_/A _2555_/Y gnd _2556_/Y vdd NAND2X1
X_2487_ _2485_/Y _2486_/Y gnd _2493_/B vdd NOR2X1
X_2625_ _2617_/Y _2619_/Y _2625_/C gnd _2625_/Y vdd AOI21X1
X_4226_ _4226_/A _4226_/B _4247_/C _4223_/Y gnd _4226_/Y vdd OAI22X1
X_3108_ _3108_/A _3108_/B gnd _3120_/B vdd NOR2X1
X_4088_ _4360_/Q _4088_/B gnd _4090_/B vdd NOR2X1
X_4157_ _4276_/A _4157_/B _4098_/S gnd _4160_/D vdd MUX2X1
X_3039_ _3143_/A gnd gnd _3143_/D gnd _3040_/C vdd AOI22X1
XFILL70960x40100 gnd vdd FILL
XSFILL29360x24100 gnd vdd FILL
XSFILL14640x44100 gnd vdd FILL
X_3390_ _3389_/Y _3390_/B gnd _3390_/Y vdd NOR2X1
X_2410_ _2307_/A _2190_/A gnd _2410_/Y vdd NAND2X1
X_2341_ _2406_/A _4588_/B gnd _3017_/A vdd OR2X2
X_4011_ _4010_/Y _4011_/B _4010_/C _4008_/Y gnd _4011_/Y vdd OAI22X1
X_2272_ _2272_/A _2272_/B gnd _2272_/Y vdd AND2X2
X_3726_ _3726_/A _3726_/B _3726_/C gnd _3726_/Y vdd OAI21X1
X_3657_ _3447_/Y gnd _3811_/A vdd INVX4
X_2539_ _2535_/Y _2539_/B _2539_/C gnd _2539_/Y vdd AOI21X1
X_2608_ _2600_/Y _2607_/Y gnd _2635_/B vdd NOR2X1
X_3588_ _3588_/A _3586_/Y _3582_/C gnd _3639_/D vdd AOI21X1
X_4209_ _4031_/A _4231_/B gnd _4209_/Y vdd NOR2X1
XSFILL44400x22100 gnd vdd FILL
XFILL71120x24100 gnd vdd FILL
X_2890_ _2890_/A _2889_/Y gnd _2890_/Y vdd NAND2X1
X_4560_ _4560_/A _4560_/B _4559_/Y gnd _4560_/Y vdd OAI21X1
X_4491_ _4489_/Y _4491_/B _4557_/C gnd _4491_/Y vdd AOI21X1
X_3511_ _3532_/A _4617_/A gnd _3517_/A vdd NAND2X1
X_2324_ _4039_/A _4217_/A gnd _2324_/Y vdd NOR2X1
X_3373_ _3372_/Y _3373_/B gnd _3374_/C vdd AND2X2
X_3442_ _3042_/Y gnd _3442_/Y vdd INVX1
XSFILL43760x50100 gnd vdd FILL
X_2255_ _2255_/A _2221_/B _2254_/Y gnd _2255_/Y vdd OAI21X1
X_2186_ _2185_/A gnd _2188_/B vdd INVX1
X_3709_ _3843_/A _3737_/B _3708_/Y gnd _3709_/Y vdd OAI21X1
X_2873_ _2874_/A _2871_/Y _2875_/B _2875_/A gnd _2922_/C vdd OAI22X1
X_3991_ _3854_/A _3943_/B gnd _3993_/B vdd NOR2X1
XSFILL14320x16100 gnd vdd FILL
X_2942_ _2965_/B _2941_/Y gnd _2982_/B vdd NAND2X1
X_4543_ _4548_/B _4541_/Y _4542_/Y gnd _4543_/Y vdd OAI21X1
X_4612_ _4612_/A _4206_/A gnd _4613_/C vdd NAND2X1
X_4474_ _4565_/Q _4470_/C _4476_/C gnd _4486_/B vdd NAND3X1
X_2238_ _2238_/A _2236_/Y gnd _3241_/A vdd NOR2X1
X_3356_ gnd gnd _3356_/Y vdd INVX1
X_3287_ gnd gnd _3287_/Y vdd INVX1
X_2307_ _2307_/A _4597_/B gnd _2307_/Y vdd AND2X2
X_3425_ _2986_/A _2986_/B gnd _3513_/B vdd OR2X2
X_2169_ _2298_/B _2298_/A gnd _2171_/B vdd AND2X2
XSFILL14640x52100 gnd vdd FILL
X_4190_ _4417_/Q _4190_/B _4199_/B gnd _4193_/D vdd MUX2X1
X_3210_ gnd _3340_/B gnd _3210_/Y vdd NAND2X1
X_3141_ _2361_/Y _3141_/B gnd _3141_/Y vdd NAND2X1
X_3072_ _2461_/Y gnd _3072_/Y vdd INVX1
X_2925_ _2925_/A _2925_/B _2924_/Y gnd _2925_/Y vdd OAI21X1
X_2856_ _2856_/A gnd _2924_/C vdd INVX1
XSFILL59440x28100 gnd vdd FILL
XBUFX2_insert19 _3564_/Y gnd _3605_/B vdd BUFX2
X_3974_ _3974_/A _4152_/B _3973_/Y gnd _4445_/D vdd AOI21X1
X_2787_ _2786_/Y _2784_/Y gnd _2787_/Y vdd NOR2X1
X_4526_ _4574_/Q _4575_/Q _4525_/Y gnd _4540_/C vdd NAND3X1
X_4457_ _4565_/Q gnd _4460_/A vdd INVX1
X_3408_ _3401_/A gnd _2113_/A vdd INVX1
XSFILL44720x48100 gnd vdd FILL
X_3339_ gnd gnd _3341_/A vdd INVX1
X_4388_ _4041_/B _4436_/CLK _4388_/D gnd vdd DFFPOSX1
XSFILL59120x10100 gnd vdd FILL
XBUFX2_insert229 _4449_/Q gnd _2786_/A vdd BUFX2
XBUFX2_insert207 _3641_/Q gnd _4124_/S vdd BUFX2
XBUFX2_insert218 _3651_/Y gnd _3671_/B vdd BUFX2
XSFILL44400x30100 gnd vdd FILL
XSFILL28880x20100 gnd vdd FILL
X_3690_ _3524_/Y gnd _3692_/A vdd INVX4
XSFILL58960x6100 gnd vdd FILL
X_2710_ _2706_/Y _2756_/B gnd _2710_/Y vdd NAND2X1
X_4311_ _3870_/A _4417_/CLK _4311_/D gnd vdd DFFPOSX1
X_2641_ _2641_/A _2637_/Y _2641_/C gnd _2641_/Y vdd NAND3X1
X_2572_ _2572_/A _2571_/A gnd _2573_/B vdd NAND2X1
X_4242_ _4064_/A _4231_/B gnd _4242_/Y vdd NOR2X1
X_4173_ _2136_/B _3951_/B _3951_/C gnd _4173_/Y vdd OAI21X1
X_3124_ _2476_/Y gnd _3124_/Y vdd INVX1
X_3055_ _3053_/Y _3341_/B _3055_/C gnd _3056_/B vdd OAI21X1
X_3957_ _4412_/Q _4135_/B _3968_/S gnd _3960_/D vdd MUX2X1
X_2839_ _2713_/A gnd _2842_/A vdd INVX1
X_2908_ _2895_/A _2898_/Y gnd _2911_/C vdd NOR2X1
X_3888_ _3788_/A _3873_/B _3888_/C gnd _4335_/D vdd AOI21X1
X_4509_ _4548_/C _4509_/B _4520_/B gnd _4511_/A vdd NAND3X1
X_3811_ _3811_/A _3823_/B _3811_/C gnd _3811_/Y vdd AOI21X1
X_3742_ _3843_/A _3740_/B _3741_/Y gnd _3742_/Y vdd OAI21X1
X_2624_ _2752_/A _2616_/Y gnd _2625_/C vdd NOR2X1
X_3673_ _3673_/A _3671_/B gnd _3673_/Y vdd NOR2X1
X_2555_ _2102_/A gnd _2555_/Y vdd INVX1
X_4225_ _3897_/A _4245_/S _4247_/C gnd _4226_/A vdd OAI21X1
X_2486_ _2475_/Y _2482_/Y gnd _2486_/Y vdd NAND2X1
X_4087_ _4124_/S gnd _4087_/Y vdd INVX8
X_3107_ _3107_/A _3341_/B _3107_/C gnd _3108_/B vdd OAI21X1
X_4156_ _4155_/Y _4156_/B _4101_/C _4153_/Y gnd _4161_/B vdd OAI22X1
X_3038_ gnd _3240_/B _3246_/C gnd _3040_/A vdd NAND3X1
XSFILL29360x40100 gnd vdd FILL
X_2271_ _2572_/A _2102_/A gnd _2272_/A vdd OR2X2
X_2340_ _2295_/A _2295_/B gnd _2991_/A vdd OR2X2
X_4010_ _4010_/A _4012_/S _4010_/C gnd _4010_/Y vdd OAI21X1
X_3725_ _4283_/A _3737_/B _3725_/C gnd _4369_/D vdd OAI21X1
XSFILL59440x36100 gnd vdd FILL
X_3656_ _3843_/A _3658_/B _3656_/C gnd _3656_/Y vdd AOI21X1
X_3587_ _3771_/A _3590_/B gnd _3588_/A vdd NAND2X1
X_2607_ _2607_/A _2606_/Y gnd _2607_/Y vdd NAND2X1
X_4208_ _4208_/A _4208_/B _4241_/S gnd _4211_/D vdd MUX2X1
X_2538_ _2538_/A _2538_/B gnd _2539_/C vdd NAND2X1
X_2469_ _2488_/A _2488_/B gnd _2472_/C vdd NAND2X1
XSFILL14800x20100 gnd vdd FILL
X_4139_ _4139_/A _4139_/B _4205_/S gnd _4141_/A vdd MUX2X1
XFILL71120x40100 gnd vdd FILL
X_4490_ _4558_/B _4595_/Y _4488_/B _4556_/D gnd _4491_/B vdd AOI22X1
X_3441_ _3518_/A _3441_/B gnd _3441_/Y vdd NAND2X1
X_3510_ _3504_/Y _3509_/Y gnd _3510_/Y vdd NAND2X1
X_2254_ _2254_/A _2229_/Y _2253_/Y gnd _2254_/Y vdd AOI21X1
X_2323_ _2321_/Y _2323_/B gnd _2323_/Y vdd NOR2X1
X_3372_ gnd _3372_/B _3372_/C gnd _3372_/Y vdd NAND3X1
X_2185_ _2185_/A _2185_/B gnd _3085_/A vdd XNOR2X1
X_3639_ _3771_/A _4300_/CLK _3639_/D gnd vdd DFFPOSX1
X_3708_ _3703_/B _3726_/B _3921_/A gnd _3708_/Y vdd OAI21X1
XFILL70960x46100 gnd vdd FILL
X_3990_ _4415_/Q _3673_/A _3992_/B gnd _3993_/D vdd MUX2X1
X_2872_ _2110_/A gnd _2875_/B vdd INVX1
X_4611_ _4611_/A gnd _4611_/Y vdd INVX1
X_2941_ _2965_/A gnd _2941_/Y vdd INVX1
X_4542_ _4558_/B _4542_/B _2150_/A _4556_/D gnd _4542_/Y vdd AOI22X1
XSFILL14320x32100 gnd vdd FILL
X_4473_ _4460_/A _4466_/Y _4479_/A gnd _4475_/C vdd OAI21X1
X_3424_ _3424_/A gnd _3427_/C vdd INVX1
X_2237_ _2235_/Y _2232_/Y gnd _2238_/A vdd NOR2X1
X_3355_ _3355_/A gnd _3357_/A vdd INVX1
X_3286_ _3286_/A _3130_/B _3285_/Y _3130_/D gnd _3290_/A vdd OAI22X1
X_2306_ _2307_/A _4597_/B gnd _2306_/Y vdd NOR2X1
X_2099_ _2779_/B gnd data_out[11] vdd BUFX2
X_2168_ _2167_/B _2168_/B _2164_/A gnd _2168_/Y vdd OAI21X1
XSFILL44400x28100 gnd vdd FILL
XSFILL29840x26100 gnd vdd FILL
X_3071_ _3069_/Y _2950_/B _3071_/C _3201_/D gnd _3071_/Y vdd OAI22X1
X_3140_ _3140_/A _3140_/B _3139_/Y gnd _3140_/Y vdd NAND3X1
X_3973_ _2190_/B _4152_/B _3649_/A gnd _3973_/Y vdd OAI21X1
X_2786_ _2786_/A _2830_/A _2786_/C _2786_/D gnd _2786_/Y vdd OAI22X1
X_2855_ _2925_/A _2925_/B _2100_/A _2854_/Y gnd _2855_/Y vdd AOI22X1
XSFILL59440x44100 gnd vdd FILL
X_2924_ _2772_/B _2859_/B _2924_/C _2745_/A gnd _2924_/Y vdd OAI22X1
X_4525_ _4506_/C _4513_/C _4513_/B gnd _4525_/Y vdd NOR3X1
X_4387_ _4208_/B _4373_/CLK _3829_/Y gnd vdd DFFPOSX1
X_3338_ _3336_/Y _3130_/B _3338_/C _3130_/D gnd _3338_/Y vdd OAI22X1
X_4456_ _4228_/C gnd _4557_/C vdd INVX4
X_3407_ _3649_/A gnd _3417_/D vdd INVX1
X_3269_ _3268_/Y _3269_/B gnd _3269_/Y vdd AND2X2
XBUFX2_insert219 _3651_/Y gnd _3658_/B vdd BUFX2
XBUFX2_insert208 _3641_/Q gnd _4166_/B vdd BUFX2
X_2640_ _2640_/A _2862_/A _2318_/B _2584_/Y gnd _2641_/C vdd AOI22X1
X_2571_ _2571_/A _2571_/B gnd _2573_/A vdd OR2X2
X_4241_ _4241_/A _4390_/Q _4241_/S gnd _4244_/D vdd MUX2X1
X_4310_ _4246_/A _4298_/CLK _3869_/Y gnd vdd DFFPOSX1
X_4172_ _4171_/Y _4172_/B _4205_/S gnd _4174_/A vdd MUX2X1
X_3123_ _3121_/Y _2950_/B _3122_/Y _3201_/D gnd _3127_/B vdd OAI22X1
X_3054_ gnd _3340_/B gnd _3055_/C vdd NAND2X1
XSFILL59760x2100 gnd vdd FILL
X_2907_ _2907_/A _2906_/Y _2903_/Y gnd _2907_/Y vdd AOI21X1
X_3956_ _3955_/Y _3956_/B _3988_/C _3953_/Y gnd _3961_/B vdd OAI22X1
X_2769_ _2832_/A _2101_/A _2100_/A _2769_/D gnd _2769_/Y vdd AOI22X1
X_4508_ _4508_/A gnd _4520_/B vdd INVX1
X_2838_ _2838_/A gnd _2838_/Y vdd INVX1
X_3887_ _3992_/A _3873_/B gnd _3888_/C vdd NOR2X1
X_4439_ _4439_/Q _4451_/CLK _4439_/D gnd vdd DFFPOSX1
XSFILL59920x40100 gnd vdd FILL
XSFILL29360x38100 gnd vdd FILL
X_3810_ _4378_/Q _3823_/B gnd _3811_/C vdd NOR2X1
X_3741_ _4313_/Q _3740_/B gnd _3741_/Y vdd NAND2X1
XSFILL29040x20100 gnd vdd FILL
X_2554_ _2554_/A _2553_/Y gnd _3332_/A vdd XNOR2X1
X_2623_ _2622_/Y _2635_/B gnd _2623_/Y vdd AND2X2
X_3672_ _3482_/Y gnd _3788_/A vdd INVX4
XSFILL14320x40100 gnd vdd FILL
X_4224_ _4046_/A _4180_/B gnd _4226_/B vdd NOR2X1
X_2485_ _2464_/A _2485_/B gnd _2485_/Y vdd NAND2X1
X_4155_ _3751_/A _4098_/S _4155_/C gnd _4155_/Y vdd OAI21X1
X_3106_ gnd _3340_/B gnd _3107_/C vdd NAND2X1
X_4086_ _3773_/A _4376_/Q _4153_/S gnd _4090_/D vdd MUX2X1
X_3037_ _2357_/Y _3141_/B gnd _3037_/Y vdd NAND2X1
X_3939_ _3939_/A _3939_/B _4027_/S gnd _3941_/A vdd MUX2X1
XSFILL58800x6100 gnd vdd FILL
XSFILL59120x16100 gnd vdd FILL
XSFILL29680x6100 gnd vdd FILL
X_2270_ _2572_/A _2102_/A gnd _2272_/B vdd NAND2X1
XSFILL29840x34100 gnd vdd FILL
X_3724_ _3726_/A _3726_/B _4187_/A gnd _3725_/C vdd OAI21X1
XSFILL59440x52100 gnd vdd FILL
X_3655_ _4393_/Q _3658_/B gnd _3656_/C vdd NOR2X1
X_3586_ _3589_/A data_in[10] gnd _3586_/Y vdd NAND2X1
X_2606_ _2604_/Y _2488_/A _2606_/C _2606_/D gnd _2606_/Y vdd AOI22X1
X_2537_ _2537_/A _2537_/B gnd _2538_/A vdd NOR2X1
X_4207_ _4207_/A _4207_/B _4206_/Y gnd _4434_/D vdd AOI21X1
X_2399_ _2399_/A _2399_/B _2396_/Y gnd _2400_/C vdd NOR3X1
X_2468_ _2633_/B gnd _2488_/B vdd INVX1
X_4138_ _4138_/A _4136_/Y _4170_/C _4138_/D gnd _4139_/A vdd OAI22X1
X_4069_ _4069_/A _4012_/S _4010_/C gnd _4070_/A vdd OAI21X1
XSFILL59600x12100 gnd vdd FILL
X_3371_ _3371_/A _2961_/A _3267_/C gnd _3373_/B vdd NAND3X1
X_3440_ _3434_/Y _3439_/Y gnd _3440_/Y vdd NAND2X1
X_2253_ _2253_/A _2253_/B _2253_/C gnd _2253_/Y vdd OAI21X1
X_2322_ _2515_/A _2516_/A gnd _2323_/B vdd AND2X2
X_2184_ _2188_/C _2184_/B gnd _2185_/B vdd NAND2X1
X_3707_ _3740_/A _3737_/B _3706_/Y gnd _3707_/Y vdd OAI21X1
X_3638_ _3702_/A _4383_/CLK _3585_/Y gnd vdd DFFPOSX1
X_3569_ _3575_/A data_in[3] gnd _3613_/B vdd NAND2X1
XSFILL59600x100 gnd vdd FILL
XSFILL29360x46100 gnd vdd FILL
X_2940_ gnd gnd _2950_/C vdd INVX1
X_2871_ _2922_/B gnd _2871_/Y vdd INVX1
X_4541_ _2150_/A _4537_/A _4548_/C gnd _4541_/Y vdd OAI21X1
X_4610_ _4621_/A _4608_/Y _4610_/C gnd _4610_/Y vdd OAI21X1
X_3354_ _3354_/A _3354_/B _3353_/Y gnd _3526_/A vdd NAND3X1
X_4472_ _4476_/C gnd _4479_/A vdd INVX1
X_3423_ _3434_/A gnd _3495_/A vdd INVX4
X_2236_ _2232_/Y _2235_/Y gnd _2236_/Y vdd AND2X2
X_3285_ gnd gnd _3285_/Y vdd INVX1
X_2305_ _2303_/Y _2304_/Y gnd _2305_/Y vdd NOR2X1
X_2167_ _2166_/Y _2167_/B gnd _2167_/Y vdd XNOR2X1
X_2098_ _2098_/A gnd data_out[10] vdd BUFX2
XSFILL59120x24100 gnd vdd FILL
XSFILL44400x44100 gnd vdd FILL
XFILL71120x46100 gnd vdd FILL
XSFILL29840x42100 gnd vdd FILL
X_3070_ gnd gnd _3071_/C vdd INVX1
X_2923_ _2864_/Y _2923_/B _2923_/C _2870_/A gnd _2929_/B vdd OAI22X1
X_3972_ _3972_/A _3972_/B _4027_/S gnd _3974_/A vdd MUX2X1
X_2785_ _2874_/A gnd _2830_/A vdd INVX1
X_2854_ _2768_/A gnd _2854_/Y vdd INVX1
X_4524_ _4522_/Y _4524_/B _4557_/C gnd _4574_/D vdd AOI21X1
X_4386_ _3826_/A _4359_/CLK _4386_/D gnd vdd DFFPOSX1
X_4455_ _4455_/Q _4451_/CLK _4084_/Y gnd vdd DFFPOSX1
X_3337_ gnd gnd _3338_/C vdd INVX1
X_3406_ _3400_/C _3406_/B _3405_/Y gnd _4462_/A vdd OAI21X1
X_2219_ _2218_/Y _2219_/B gnd _2219_/Y vdd NOR2X1
X_3199_ _3199_/A gnd _3201_/A vdd INVX1
X_3268_ gnd _3346_/B _3268_/C gnd _3268_/Y vdd NAND3X1
XBUFX2_insert209 _3641_/Q gnd _4252_/S vdd BUFX2
XSFILL59600x20100 gnd vdd FILL
X_2570_ _2661_/A gnd _2571_/A vdd INVX1
X_4240_ _4238_/Y _4240_/B _4239_/Y gnd _4240_/Y vdd AOI21X1
X_4171_ _4170_/Y _4171_/B _4170_/C _4171_/D gnd _4171_/Y vdd OAI22X1
X_3122_ gnd gnd _3122_/Y vdd INVX1
XSFILL14320x38100 gnd vdd FILL
X_3053_ gnd gnd _3053_/Y vdd INVX1
X_2906_ _2906_/A _2906_/B gnd _2906_/Y vdd NAND2X1
X_3955_ _4133_/A _3968_/S _3988_/C gnd _3955_/Y vdd OAI21X1
X_3886_ _3752_/A _3879_/B _3885_/Y gnd _3886_/Y vdd AOI21X1
X_2768_ _2768_/A gnd _2769_/D vdd INVX1
X_2837_ _2837_/A _2837_/B _2837_/C gnd _2844_/C vdd AOI21X1
X_4438_ _4438_/Q _4451_/CLK _4438_/D gnd vdd DFFPOSX1
X_4507_ _4506_/C _4513_/B gnd _4508_/A vdd NOR2X1
X_2699_ _2890_/A _2699_/B gnd _2699_/Y vdd NAND2X1
X_4369_ _4187_/A _4417_/CLK _4369_/D gnd vdd DFFPOSX1
X_3740_ _3740_/A _3740_/B _3739_/Y gnd _4312_/D vdd OAI21X1
X_2553_ _2572_/A _2102_/A gnd _2553_/Y vdd XNOR2X1
X_2622_ _2620_/Y _2621_/Y _2622_/C gnd _2622_/Y vdd NOR3X1
X_3671_ _3752_/A _3671_/B _3670_/Y gnd _4398_/D vdd AOI21X1
X_4223_ _4045_/A _3688_/A _4245_/S gnd _4223_/Y vdd MUX2X1
X_3105_ gnd gnd _3107_/A vdd INVX1
X_4085_ _4085_/A gnd _4205_/S vdd INVX8
X_2484_ _2488_/A _2633_/B gnd _2485_/B vdd XNOR2X1
X_4154_ _4366_/Q _4158_/B gnd _4156_/B vdd NOR2X1
X_3036_ _3031_/Y _3036_/B _3036_/C gnd _3036_/Y vdd NAND3X1
X_3869_ _3902_/A _3862_/B _3869_/C gnd _3869_/Y vdd OAI21X1
XSFILL14800x34100 gnd vdd FILL
X_3938_ _3938_/A _3936_/Y _3934_/C _3935_/Y gnd _3939_/A vdd OAI22X1
XSFILL44400x52100 gnd vdd FILL
XSFILL59600x2100 gnd vdd FILL
XSFILL29840x50100 gnd vdd FILL
X_3723_ _4281_/A _3737_/B _3723_/C gnd _4368_/D vdd OAI21X1
X_3654_ _3440_/Y gnd _3843_/A vdd INVX4
X_3585_ _3585_/A _3583_/Y _3582_/C gnd _3585_/Y vdd AOI21X1
X_2467_ _2633_/B _2466_/Y gnd _2474_/A vdd NAND2X1
X_2605_ _2891_/A gnd _2606_/C vdd INVX1
X_2536_ _2482_/A _2482_/B gnd _2537_/B vdd XOR2X1
XSFILL59760x8100 gnd vdd FILL
X_4206_ _4206_/A _4207_/B _4206_/C gnd _4206_/Y vdd OAI21X1
X_4068_ _4246_/A _4020_/B gnd _4068_/Y vdd NOR2X1
X_2398_ _2421_/A _4184_/A gnd _2399_/B vdd XOR2X1
X_4137_ _3881_/A _4166_/B _4170_/C gnd _4138_/A vdd OAI21X1
XSFILL44880x24100 gnd vdd FILL
XSFILL29360x100 gnd vdd FILL
X_3019_ _3019_/A _2950_/B _3018_/Y _3201_/D gnd _3023_/B vdd OAI22X1
XSFILL59920x46100 gnd vdd FILL
X_3370_ _3370_/A _3267_/C _3292_/C gnd _3374_/B vdd NAND3X1
X_2321_ _2515_/A _2516_/A gnd _2321_/Y vdd NOR2X1
X_2252_ _2252_/A _2252_/B _2233_/Y gnd _2253_/C vdd OAI21X1
X_2183_ _2187_/A _2193_/B gnd _2184_/B vdd OR2X2
XSFILL14320x46100 gnd vdd FILL
XSFILL29520x6100 gnd vdd FILL
X_3637_ _2965_/A _3632_/CLK _3637_/D gnd vdd DFFPOSX1
X_3706_ _3706_/A _3726_/B _4360_/Q gnd _3706_/Y vdd OAI21X1
X_2519_ _2252_/A _2520_/A gnd _2519_/Y vdd NOR2X1
X_3568_ _3982_/C _3574_/B gnd _3570_/A vdd NAND2X1
X_3499_ _3513_/A _3513_/B _3499_/C gnd _3499_/Y vdd OAI21X1
XSFILL44880x6100 gnd vdd FILL
X_2870_ _2870_/A gnd _2878_/A vdd INVX1
X_4540_ _4540_/A _4540_/B _4540_/C gnd _4548_/B vdd NOR3X1
X_4471_ _4471_/A _4469_/Y _4557_/C gnd _4566_/D vdd AOI21X1
X_3353_ _3353_/A _3352_/Y gnd _3353_/Y vdd NOR2X1
X_3284_ gnd gnd _3286_/A vdd INVX1
X_2304_ _2193_/B _2187_/A gnd _2304_/Y vdd AND2X2
X_3422_ _3422_/A _3422_/B gnd _3422_/Y vdd NAND2X1
X_2235_ _2235_/A _2233_/Y gnd _2235_/Y vdd NOR2X1
X_2097_ _2442_/A gnd data_out[1] vdd BUFX2
X_2166_ _2168_/B _2164_/Y gnd _2166_/Y vdd NOR2X1
XSFILL29520x22100 gnd vdd FILL
X_2999_ gnd gnd _3000_/C vdd INVX1
XSFILL14800x42100 gnd vdd FILL
XFILL70960x100 gnd vdd FILL
XSFILL59600x18100 gnd vdd FILL
X_2922_ _2922_/A _2922_/B _2922_/C gnd _2923_/C vdd OAI21X1
X_2853_ _2772_/B gnd _2925_/A vdd INVX1
X_3971_ _3970_/Y _3969_/Y _3988_/C _3971_/D gnd _3972_/A vdd OAI22X1
X_2784_ _2874_/A _2784_/B _2783_/Y gnd _2784_/Y vdd OAI21X1
X_4454_ _4454_/Q _4451_/CLK _4073_/Y gnd vdd DFFPOSX1
X_4523_ _4558_/B _4610_/Y _4574_/Q _4556_/D gnd _4524_/B vdd AOI22X1
X_4385_ _4186_/B _4417_/CLK _3825_/Y gnd vdd DFFPOSX1
X_3267_ _3267_/A _3345_/B _3267_/C gnd _3269_/B vdd NAND3X1
X_3336_ gnd gnd _3336_/Y vdd INVX1
X_3405_ _3405_/A _3400_/C _3413_/A gnd _3405_/Y vdd AOI21X1
X_2149_ _2158_/A _2147_/Y _2148_/Y gnd _2149_/Y vdd OAI21X1
X_2218_ _2782_/A _2218_/B gnd _2218_/Y vdd NOR2X1
X_3198_ _3198_/A _3198_/B _3197_/Y gnd _3484_/A vdd NAND3X1
X_4170_ _3992_/A _4166_/B _4170_/C gnd _4170_/Y vdd OAI21X1
X_3121_ _3121_/A gnd _3121_/Y vdd INVX1
X_3052_ _3050_/Y _3130_/B _3052_/C _3130_/D gnd _3056_/A vdd OAI22X1
X_2836_ _2769_/Y _2836_/B _2836_/C gnd _2837_/C vdd OAI21X1
X_2905_ _2619_/A _2905_/B gnd _2907_/A vdd NAND2X1
X_3954_ _3714_/C _3943_/B gnd _3956_/B vdd NOR2X1
X_3885_ _4334_/Q _3879_/B gnd _3885_/Y vdd NOR2X1
X_4437_ _4437_/Q _4417_/CLK _4240_/Y gnd vdd DFFPOSX1
X_2767_ _2772_/B gnd _2832_/A vdd INVX1
X_4506_ _4499_/Y _4495_/Y _4506_/C gnd _4509_/B vdd OAI21X1
X_2698_ _2723_/B gnd _2699_/B vdd INVX1
X_4368_ _4176_/A _4373_/CLK _4368_/D gnd vdd DFFPOSX1
X_3319_ _3319_/A _2961_/A _3267_/C gnd _3321_/B vdd NAND3X1
X_4299_ _3947_/A _4298_/CLK _3847_/Y gnd vdd DFFPOSX1
XSFILL29840x48100 gnd vdd FILL
X_3670_ _4157_/B _3658_/B gnd _3670_/Y vdd NOR2X1
X_4222_ _4222_/A _4222_/B _4247_/C _4219_/Y gnd _4227_/B vdd OAI22X1
X_2552_ _2529_/Y _2552_/B _2551_/Y gnd _2554_/A vdd AOI21X1
X_2621_ _2752_/A _2616_/Y _2619_/A _2618_/Y gnd _2621_/Y vdd OAI22X1
X_2483_ _2481_/Y _2482_/Y gnd _2483_/Y vdd XNOR2X1
X_4084_ _4084_/A _4207_/B _4083_/Y gnd _4084_/Y vdd AOI21X1
X_3104_ _3102_/Y _3130_/B _3104_/C _3130_/D gnd _3108_/A vdd OAI22X1
X_4153_ _4153_/A _4153_/B _4153_/S gnd _4153_/Y vdd MUX2X1
X_3035_ _3035_/A _3033_/Y gnd _3036_/C vdd AND2X2
X_3937_ _3877_/A _4030_/S _3934_/C gnd _3938_/A vdd OAI21X1
XSFILL29520x30100 gnd vdd FILL
X_3799_ _3799_/A _3803_/B gnd _3800_/C vdd NAND2X1
X_3868_ _4246_/A _3862_/B gnd _3869_/C vdd NAND2X1
X_2819_ _2633_/B _2817_/A gnd _2823_/A vdd NOR2X1
X_3722_ _3732_/A _3726_/B _4176_/A gnd _3723_/C vdd OAI21X1
X_2604_ _2723_/B gnd _2604_/Y vdd INVX1
X_3653_ _3740_/A _3658_/B _3653_/C gnd _3653_/Y vdd AOI21X1
X_4205_ _4204_/Y _4205_/B _4205_/S gnd _4207_/A vdd MUX2X1
X_2535_ _2445_/B _2452_/Y _2535_/C gnd _2535_/Y vdd NAND3X1
X_3584_ _3702_/A _3590_/B gnd _3585_/A vdd NAND2X1
X_2466_ _2488_/A gnd _2466_/Y vdd INVX1
X_4067_ _4292_/A _4245_/B _4012_/S gnd _4070_/D vdd MUX2X1
X_2397_ _4050_/A _2351_/B gnd _2399_/A vdd XOR2X1
X_4136_ _4300_/Q _4088_/B gnd _4136_/Y vdd NOR2X1
X_3018_ gnd gnd _3018_/Y vdd INVX1
XSFILL14000x26100 gnd vdd FILL
X_2320_ _2320_/A _2320_/B gnd _3214_/A vdd NOR2X1
X_2251_ _2251_/A gnd _2254_/A vdd INVX1
X_2182_ _2187_/A _2193_/B gnd _2188_/C vdd NAND2X1
X_3567_ _3565_/Y _3611_/B _3582_/C gnd _3567_/Y vdd AOI21X1
X_3636_ _2965_/B _3632_/CLK _3636_/D gnd vdd DFFPOSX1
XBUFX2_insert190 _4426_/Q gnd _4588_/B vdd BUFX2
X_3705_ _3702_/A _3704_/A gnd _3726_/B vdd NAND2X1
X_2518_ _2252_/B gnd _2520_/A vdd INVX1
X_2449_ _2614_/C gnd _2450_/B vdd INVX1
X_3498_ _3498_/A gnd _3499_/C vdd INVX1
X_4119_ _4119_/A _4130_/B _4118_/Y gnd _4426_/D vdd AOI21X1
XSFILL59120x38100 gnd vdd FILL
XSFILL59600x8100 gnd vdd FILL
X_4470_ _4558_/B _4586_/Y _4470_/C _4556_/D gnd _4471_/A vdd AOI22X1
X_3421_ _3421_/Q _3632_/CLK _3421_/D gnd vdd DFFPOSX1
X_2234_ _2778_/A _2098_/A gnd _2235_/A vdd NOR2X1
X_3283_ _3283_/A _3283_/B gnd _3302_/A vdd NOR2X1
X_3352_ _3352_/A _3352_/B _3351_/Y gnd _3352_/Y vdd NAND3X1
X_2303_ _2193_/B _2187_/A gnd _2303_/Y vdd NOR2X1
X_2096_ _2794_/A gnd data_out[0] vdd BUFX2
XSFILL59280x8100 gnd vdd FILL
X_2165_ _2392_/B _2295_/A gnd _2168_/B vdd NOR2X1
X_2998_ gnd gnd _2998_/Y vdd INVX1
X_3619_ _3618_/Y _3579_/B _3579_/C gnd _3632_/D vdd AOI21X1
X_4599_ _3469_/B gnd _4601_/B vdd INVX1
XSFILL43920x46100 gnd vdd FILL
X_3970_ _3970_/A _3968_/S _3988_/C gnd _3970_/Y vdd OAI21X1
X_2921_ _2829_/B _2921_/B gnd _2923_/B vdd NOR2X1
X_2783_ _2786_/C _2786_/D gnd _2783_/Y vdd NAND2X1
X_2852_ _2846_/Y _2848_/Y _2852_/C gnd _2852_/Y vdd NAND3X1
XFILL71280x14100 gnd vdd FILL
X_4453_ _4453_/Q _4451_/CLK _4453_/D gnd vdd DFFPOSX1
X_4384_ _3997_/B _4373_/CLK _3823_/Y gnd vdd DFFPOSX1
X_4522_ _4528_/A _4528_/B _4521_/Y gnd _4522_/Y vdd OAI21X1
X_3404_ _3396_/B _2965_/B _3384_/A gnd _3405_/A vdd NAND3X1
X_2217_ _2216_/Y gnd _2219_/B vdd INVX1
X_3335_ _3334_/Y _3335_/B gnd _3354_/A vdd NOR2X1
X_3266_ _3266_/A _3188_/B _3188_/C gnd _3270_/B vdd NAND3X1
X_3197_ _3197_/A _3196_/Y gnd _3197_/Y vdd NOR2X1
XSFILL44720x6100 gnd vdd FILL
X_2148_ _2158_/A _2374_/B gnd _2148_/Y vdd NAND2X1
X_3120_ _3101_/Y _3120_/B _3120_/C gnd _3463_/A vdd NAND3X1
X_3051_ gnd gnd _3052_/C vdd INVX1
X_3953_ _4131_/A _3814_/A _3968_/S gnd _3953_/Y vdd MUX2X1
X_2766_ _2766_/A _2766_/B gnd _2766_/Y vdd NOR2X1
X_2835_ _2849_/A _2765_/B _2835_/C gnd _2836_/C vdd AOI21X1
XSFILL29520x28100 gnd vdd FILL
X_2904_ _2794_/A gnd _2905_/B vdd INVX1
X_3884_ _3717_/A _3873_/B _3884_/C gnd _3884_/Y vdd AOI21X1
XSFILL30000x16100 gnd vdd FILL
X_4436_ _4436_/Q _4436_/CLK _4229_/Y gnd vdd DFFPOSX1
X_4505_ _2135_/A gnd _4506_/C vdd INVX2
X_3318_ _3318_/A _3267_/C _3292_/C gnd _3322_/B vdd NAND3X1
X_2697_ _2723_/A _2723_/B _2891_/A _2696_/Y gnd _2702_/C vdd AOI22X1
X_4367_ _4367_/Q _4383_/CLK _3721_/Y gnd vdd DFFPOSX1
XSFILL14800x48100 gnd vdd FILL
X_4298_ _3936_/A _4298_/CLK _4298_/D gnd vdd DFFPOSX1
X_3249_ _3249_/A _3248_/Y gnd _3250_/C vdd NOR2X1
XSFILL14160x4100 gnd vdd FILL
XSFILL29200x10100 gnd vdd FILL
X_2620_ _2617_/Y _2619_/Y gnd _2620_/Y vdd NAND2X1
X_4221_ _4221_/A _4245_/S _4247_/C gnd _4222_/A vdd OAI21X1
X_2551_ _2545_/Y _2532_/Y _2547_/Y gnd _2551_/Y vdd OAI21X1
X_2482_ _2482_/A _2482_/B gnd _2482_/Y vdd XNOR2X1
X_4083_ _2849_/A _4207_/B _4206_/C gnd _4083_/Y vdd OAI21X1
X_3103_ gnd gnd _3104_/C vdd INVX1
X_4152_ _4152_/A _4152_/B _4151_/Y gnd _4429_/D vdd AOI21X1
X_3034_ gnd _3372_/B _3372_/C gnd _3035_/A vdd NAND3X1
X_3936_ _3936_/A _3932_/B gnd _3936_/Y vdd NOR2X1
X_2749_ _2678_/Y _2685_/Y gnd _2750_/A vdd NAND2X1
X_3798_ _3764_/A _3792_/B _3797_/Y gnd _4356_/D vdd OAI21X1
X_3867_ _3692_/A _3866_/B _3867_/C gnd _4309_/D vdd OAI21X1
X_2818_ _2465_/B gnd _2820_/A vdd INVX1
XSFILL44880x38100 gnd vdd FILL
X_4419_ _4212_/A _4298_/CLK _4419_/D gnd vdd DFFPOSX1
XSFILL59600x42100 gnd vdd FILL
XSFILL44560x20100 gnd vdd FILL
X_2534_ _2529_/Y _2533_/Y gnd _3280_/A vdd XNOR2X1
X_3583_ _3589_/A data_in[9] gnd _3583_/Y vdd NAND2X1
X_2603_ _2633_/A _2723_/B _2891_/A _2603_/D gnd _2607_/A vdd AOI22X1
X_3721_ _3788_/A _3737_/B _3720_/Y gnd _3721_/Y vdd OAI21X1
X_3652_ _4392_/Q _3658_/B gnd _3653_/C vdd NOR2X1
XFILL71280x22100 gnd vdd FILL
X_4204_ _4204_/A _4202_/Y _4254_/C _4204_/D gnd _4204_/Y vdd OAI22X1
X_2465_ _2465_/A _2465_/B _2464_/Y gnd _2465_/Y vdd OAI21X1
X_4135_ _4412_/Q _4135_/B _4166_/B gnd _4138_/D vdd MUX2X1
X_2396_ _2396_/A _2392_/Y _2394_/Y _2395_/Y gnd _2396_/Y vdd OAI22X1
X_4066_ _4066_/A _4064_/Y _4065_/C _4063_/Y gnd _4071_/B vdd OAI22X1
X_3017_ _3017_/A gnd _3019_/A vdd INVX1
X_3919_ _3919_/A _3941_/B _3918_/Y gnd _4440_/D vdd AOI21X1
X_2250_ _2232_/A _2251_/A gnd _2255_/A vdd OR2X2
X_2181_ _2278_/B _2278_/A gnd _2185_/A vdd NAND2X1
X_3704_ _3704_/A _3703_/Y gnd _3737_/B vdd NAND2X1
X_2517_ _2516_/Y _2514_/B gnd _2517_/Y vdd NAND2X1
XSFILL29520x36100 gnd vdd FILL
X_3497_ _3518_/A _4611_/A gnd _3503_/A vdd NAND2X1
XBUFX2_insert180 _3625_/Q gnd _4628_/A vdd BUFX2
X_3566_ data_in[2] _3589_/A gnd _3611_/B vdd NAND2X1
X_3635_ _2986_/A _3632_/CLK _3597_/Y gnd vdd DFFPOSX1
XSFILL14480x14100 gnd vdd FILL
XBUFX2_insert191 _4426_/Q gnd _2298_/B vdd BUFX2
X_2379_ _4061_/A _4239_/A gnd _2383_/B vdd AND2X2
X_2448_ _2447_/Y _2446_/Y _2440_/A gnd _2535_/C vdd OAI21X1
X_4118_ _4588_/B _4130_/B _4162_/C gnd _4118_/Y vdd OAI21X1
X_4049_ _4048_/Y _4049_/B _4027_/S gnd _4049_/Y vdd MUX2X1
X_3351_ _3143_/A gnd gnd _3143_/D gnd _3351_/Y vdd AOI22X1
X_3420_ _3413_/A _3632_/CLK _3420_/D gnd vdd DFFPOSX1
X_2233_ _2778_/A _2098_/A gnd _2233_/Y vdd AND2X2
X_3282_ _3280_/Y _3204_/B _3281_/Y _3204_/D gnd _3283_/A vdd OAI22X1
X_2302_ _2300_/Y _2302_/B gnd _2302_/Y vdd NOR2X1
X_2164_ _2164_/A gnd _2164_/Y vdd INVX1
X_2095_ _2143_/Y gnd adrs_bus[9] vdd BUFX2
X_2997_ _2996_/Y _2997_/B gnd _2997_/Y vdd NOR2X1
X_3618_ _3561_/B _3574_/B gnd _3618_/Y vdd NAND2X1
X_3549_ _3560_/B gnd _3550_/B vdd INVX1
X_4598_ _4586_/A _4596_/Y _4597_/Y gnd _4598_/Y vdd OAI21X1
XSFILL59600x50100 gnd vdd FILL
X_2920_ _2912_/Y _2920_/B _2919_/Y gnd _2920_/Y vdd AOI21X1
X_2782_ _2782_/A gnd _2786_/D vdd INVX1
X_2851_ _2926_/B _2762_/A _2762_/C _2851_/D gnd _2852_/C vdd AOI22X1
X_4521_ _4521_/A _4548_/C gnd _4521_/Y vdd AND2X2
X_4452_ _4452_/Q _4436_/CLK _4051_/Y gnd vdd DFFPOSX1
X_3334_ _3334_/A _3204_/B _3333_/Y _3204_/D gnd _3334_/Y vdd OAI22X1
X_3403_ _3413_/A _3406_/B _3402_/Y gnd _4560_/A vdd OAI21X1
X_4383_ _3820_/A _4383_/CLK _4383_/D gnd vdd DFFPOSX1
X_2147_ _2147_/A gnd _2147_/Y vdd INVX1
X_2216_ _2782_/A _2218_/B gnd _2216_/Y vdd NAND2X1
X_3265_ gnd _3343_/B gnd _3270_/A vdd NAND2X1
X_3196_ _3194_/Y _3196_/B _3195_/Y gnd _3196_/Y vdd NAND3X1
X_3050_ gnd gnd _3050_/Y vdd INVX1
X_2903_ _2906_/A _2906_/B gnd _2903_/Y vdd NOR2X1
X_3883_ _3970_/A _3873_/B gnd _3884_/C vdd NOR2X1
X_3952_ _3952_/A _3941_/B _3951_/Y gnd _4443_/D vdd AOI21X1
X_2834_ _2762_/B _2762_/A _2833_/Y gnd _2835_/C vdd AOI21X1
X_2765_ _2849_/A _2765_/B _2764_/Y _2761_/A gnd _2766_/B vdd OAI22X1
X_4504_ _4504_/A _4504_/B _4557_/C gnd _4571_/D vdd AOI21X1
X_2696_ _2913_/D gnd _2696_/Y vdd INVX1
X_4435_ _4435_/Q _4451_/CLK _4218_/Y gnd vdd DFFPOSX1
XSFILL29520x44100 gnd vdd FILL
X_3317_ gnd _3343_/B gnd _3317_/Y vdd NAND2X1
X_4297_ _4297_/Q _4297_/CLK _4297_/D gnd vdd DFFPOSX1
X_4366_ _4366_/Q _4345_/CLK _3719_/Y gnd vdd DFFPOSX1
X_3179_ _3178_/Y _3179_/B gnd _3198_/A vdd NOR2X1
X_3248_ _3248_/A _3248_/B _3247_/Y gnd _3248_/Y vdd NAND3X1
XSFILL44080x40100 gnd vdd FILL
XSFILL44560x18100 gnd vdd FILL
X_2550_ _2533_/Y _2548_/Y gnd _2552_/B vdd NOR2X1
X_4220_ _4042_/A _4180_/B gnd _4222_/B vdd NOR2X1
X_2481_ _2491_/B _2480_/Y gnd _2481_/Y vdd NOR2X1
X_4151_ _4597_/B _4152_/B _3649_/A gnd _4151_/Y vdd OAI21X1
X_4082_ _4082_/A _4077_/Y _4027_/S gnd _4084_/A vdd MUX2X1
X_3102_ gnd gnd _3102_/Y vdd INVX1
X_3033_ _2172_/Y _3007_/B _3032_/B gnd _3033_/Y vdd NAND3X1
X_3866_ _4057_/A _3866_/B gnd _3867_/C vdd NAND2X1
X_3935_ _3935_/A _3935_/B _4030_/S gnd _3935_/Y vdd MUX2X1
X_4418_ _4418_/Q _4359_/CLK _4285_/Y gnd vdd DFFPOSX1
X_2679_ _2922_/B gnd _2679_/Y vdd INVX1
X_2748_ _2748_/A _2740_/Y _2747_/Y gnd _2748_/Y vdd NAND3X1
X_3797_ _4041_/A _3792_/B gnd _3797_/Y vdd NAND2X1
X_2817_ _2817_/A _2633_/B _2465_/B _2817_/D gnd _2817_/Y vdd AOI22X1
XSFILL60080x22100 gnd vdd FILL
X_4349_ _4142_/A _4383_/CLK _3784_/Y gnd vdd DFFPOSX1
XSFILL14000x4100 gnd vdd FILL
X_3720_ _3706_/A _3726_/B _4367_/Q gnd _3720_/Y vdd OAI21X1
X_2533_ _2533_/A _2532_/Y gnd _2533_/Y vdd NAND2X1
X_3582_ _3582_/A _3621_/B _3582_/C gnd _3582_/Y vdd AOI21X1
X_2602_ _2913_/D gnd _2603_/D vdd INVX1
X_3651_ _3651_/A _3651_/B gnd _3651_/Y vdd AND2X2
X_4203_ _4025_/A _4199_/B _4254_/C gnd _4204_/A vdd OAI21X1
X_2464_ _2464_/A _2474_/D gnd _2464_/Y vdd NAND2X1
X_4134_ _4134_/A _4132_/Y _4170_/C _4131_/Y gnd _4139_/B vdd OAI22X1
X_2395_ _2395_/A _2394_/B gnd _2395_/Y vdd NOR2X1
X_4065_ _3767_/A _4052_/S _4065_/C gnd _4066_/A vdd OAI21X1
X_3016_ _2997_/Y _3016_/B _3016_/C gnd _3435_/A vdd NAND3X1
X_3849_ _4273_/A _3852_/B _3848_/Y gnd _3849_/Y vdd OAI21X1
X_3918_ _2429_/A _3941_/B _4162_/C gnd _3918_/Y vdd OAI21X1
XSFILL45040x38100 gnd vdd FILL
X_2180_ _2179_/Y _2171_/B _2180_/C gnd _2278_/B vdd AOI21X1
XBUFX2_insert192 _4454_/Q gnd _2661_/A vdd BUFX2
X_3634_ _2986_/B _3632_/CLK _3634_/D gnd vdd DFFPOSX1
XBUFX2_insert170 _4441_/Q gnd _2295_/A vdd BUFX2
XBUFX2_insert181 _3625_/Q gnd _4586_/A vdd BUFX2
X_3703_ _3702_/Y _3703_/B gnd _3703_/Y vdd NOR2X1
X_2516_ _2516_/A _2516_/B gnd _2516_/Y vdd NAND2X1
XSFILL14480x30100 gnd vdd FILL
X_3496_ _3496_/A _3495_/Y gnd _3496_/Y vdd NAND2X1
X_3565_ _3968_/S _3590_/B gnd _3565_/Y vdd NAND2X1
X_2447_ _2906_/A _2437_/B gnd _2447_/Y vdd NOR2X1
X_4048_ _4047_/Y _4046_/Y _4004_/C _4045_/Y gnd _4048_/Y vdd OAI22X1
X_4117_ _4117_/A _4117_/B _4205_/S gnd _4119_/A vdd MUX2X1
X_2378_ _2406_/A _4588_/B gnd _2378_/Y vdd XOR2X1
XSFILL44560x26100 gnd vdd FILL
XSFILL59760x100 gnd vdd FILL
XSFILL59600x48100 gnd vdd FILL
X_3350_ gnd _3194_/B _3194_/C gnd _3352_/A vdd NAND3X1
X_2301_ _2301_/A _2301_/B gnd _2302_/B vdd AND2X2
X_2232_ _2232_/A _2221_/B _2230_/Y gnd _2232_/Y vdd OAI21X1
XSFILL43600x42100 gnd vdd FILL
X_3281_ gnd gnd _3281_/Y vdd INVX1
XFILL71280x28100 gnd vdd FILL
X_2163_ _2295_/B _2295_/A gnd _2164_/A vdd NAND2X1
X_2094_ _2140_/Y gnd adrs_bus[8] vdd BUFX2
X_3617_ _3617_/A _3576_/B _3570_/C gnd _3631_/D vdd AOI21X1
X_2996_ _2994_/Y _3204_/B _2995_/Y _3204_/D gnd _2996_/Y vdd OAI22X1
X_4597_ _3562_/A _4597_/B gnd _4597_/Y vdd NAND2X1
XSFILL60080x30100 gnd vdd FILL
X_3479_ data_in[7] gnd _3480_/A vdd INVX1
X_3548_ _3562_/A _3547_/Y gnd _4593_/A vdd NOR2X1
X_2850_ _2761_/A gnd _2851_/D vdd INVX1
X_4451_ _4451_/Q _4451_/CLK _4040_/Y gnd vdd DFFPOSX1
X_2781_ _2922_/B gnd _2784_/B vdd INVX1
X_4520_ _4513_/C _4520_/B _4528_/A gnd _4521_/A vdd OAI21X1
X_3333_ gnd gnd _3333_/Y vdd INVX1
X_3264_ _3264_/A _3263_/Y gnd _3276_/B vdd NOR2X1
X_4382_ _4153_/B _4383_/CLK _4382_/D gnd vdd DFFPOSX1
X_3402_ _3400_/C gnd _3402_/Y vdd INVX1
X_2146_ _2158_/A _2144_/Y _2145_/Y gnd _2146_/Y vdd OAI21X1
X_3195_ _3143_/A gnd gnd _3143_/D gnd _3195_/Y vdd AOI22X1
X_2215_ _2215_/A _2185_/A _2280_/A gnd _2221_/B vdd AOI21X1
X_2979_ _2979_/A _2977_/Y gnd _2980_/C vdd AND2X2
XSFILL29200x24100 gnd vdd FILL
X_2833_ _2761_/A _2764_/Y gnd _2833_/Y vdd NAND2X1
X_2902_ _2711_/A gnd _2906_/B vdd INVX1
X_3951_ _2377_/A _3951_/B _3951_/C gnd _3951_/Y vdd OAI21X1
X_3882_ _4273_/A _3873_/B _3882_/C gnd _4332_/D vdd AOI21X1
X_4434_ _4434_/Q _4451_/CLK _4434_/D gnd vdd DFFPOSX1
X_2764_ _2762_/C gnd _2764_/Y vdd INVX1
X_4503_ _4558_/B _4601_/Y _4501_/B _4556_/D gnd _4504_/B vdd AOI22X1
X_2695_ _2890_/A gnd _2723_/A vdd INVX1
X_3247_ _3143_/A gnd gnd _3143_/D gnd _3247_/Y vdd AOI22X1
X_3316_ _3312_/Y _3315_/Y gnd _3316_/Y vdd NOR2X1
X_4365_ _4365_/Q _4383_/CLK _4365_/D gnd vdd DFFPOSX1
X_4296_ _3840_/A _4297_/CLK _4296_/D gnd vdd DFFPOSX1
X_3178_ _3178_/A _3204_/B _3178_/C _3204_/D gnd _3178_/Y vdd OAI22X1
X_2129_ _4495_/A gnd _2131_/B vdd INVX1
XSFILL59280x14100 gnd vdd FILL
XSFILL44560x34100 gnd vdd FILL
X_2480_ _2537_/A _2476_/A gnd _2480_/Y vdd NOR2X1
XSFILL43600x50100 gnd vdd FILL
X_4081_ _4081_/A _4079_/Y _4021_/C _4081_/D gnd _4082_/A vdd OAI22X1
X_4150_ _4149_/Y _4150_/B _4205_/S gnd _4152_/A vdd MUX2X1
X_3101_ _3100_/Y _3101_/B gnd _3101_/Y vdd NOR2X1
XFILL71280x36100 gnd vdd FILL
X_3032_ _2299_/Y _3032_/B _2947_/A gnd _3036_/B vdd NAND3X1
X_3796_ _3729_/A _3802_/B _3796_/C gnd _3796_/Y vdd OAI21X1
X_3865_ _3764_/A _3866_/B _3865_/C gnd _4308_/D vdd OAI21X1
X_3934_ _3934_/A _3932_/Y _3934_/C _3934_/D gnd _3939_/B vdd OAI22X1
X_2816_ _2606_/D gnd _2817_/D vdd INVX1
X_4417_ _4417_/Q _4417_/CLK _4283_/Y gnd vdd DFFPOSX1
X_2678_ _2734_/C _2678_/B gnd _2678_/Y vdd NOR2X1
X_2747_ _2665_/A _2663_/Y _2746_/Y gnd _2747_/Y vdd AOI21X1
X_4348_ _4131_/A _4383_/CLK _3782_/Y gnd vdd DFFPOSX1
X_4279_ _3788_/A _4269_/B _4278_/Y gnd _4279_/Y vdd AOI21X1
XSFILL29840x2100 gnd vdd FILL
X_3650_ _3702_/A _3706_/A gnd _3651_/A vdd NOR2X1
X_4202_ _4024_/A _4198_/B gnd _4202_/Y vdd NOR2X1
X_2532_ _2530_/Y _2351_/A gnd _2532_/Y vdd OR2X2
X_3581_ _3564_/A data_in[7] gnd _3621_/B vdd NAND2X1
X_2601_ _2890_/A gnd _2633_/A vdd INVX1
X_2463_ _2606_/D _2465_/B gnd _2464_/A vdd XNOR2X1
X_4064_ _4064_/A _4002_/B gnd _4064_/Y vdd NOR2X1
X_4133_ _4133_/A _4166_/B _4170_/C gnd _4134_/A vdd OAI21X1
X_2394_ _2307_/A _2394_/B gnd _2394_/Y vdd AND2X2
X_3015_ _3015_/A _3015_/B gnd _3016_/C vdd NOR2X1
XSFILL14480x28100 gnd vdd FILL
X_3917_ _3649_/C _3916_/Y gnd _3917_/Y vdd NOR2X1
X_3848_ _4300_/Q _3852_/B gnd _3848_/Y vdd NAND2X1
X_3779_ _4347_/Q _3775_/B gnd _3780_/C vdd NAND2X1
XSFILL44080x46100 gnd vdd FILL
XSFILL29200x32100 gnd vdd FILL
XBUFX2_insert160 _4435_/Q gnd _2862_/A vdd BUFX2
XBUFX2_insert193 _4454_/Q gnd _2761_/A vdd BUFX2
XBUFX2_insert182 _3625_/Q gnd _4621_/A vdd BUFX2
X_3633_ _3553_/A _3632_/CLK _3633_/D gnd vdd DFFPOSX1
XBUFX2_insert171 _4441_/Q gnd _2711_/A vdd BUFX2
X_3702_ _3702_/A gnd _3702_/Y vdd INVX1
X_2515_ _2515_/A gnd _2516_/B vdd INVX1
X_3495_ _3495_/A _3494_/Y _3492_/Y gnd _3495_/Y vdd NAND3X1
X_3564_ _3564_/A gnd _3564_/Y vdd INVX8
X_2446_ _2434_/Y _2794_/A gnd _2446_/Y vdd AND2X2
X_4047_ _3897_/A _4036_/B _4004_/C gnd _4047_/Y vdd OAI21X1
X_4116_ _4116_/A _4116_/B _4111_/C _4113_/Y gnd _4117_/A vdd OAI22X1
X_2377_ _2377_/A _4591_/B gnd _2377_/Y vdd XOR2X1
XSFILL14960x24100 gnd vdd FILL
XFILL71280x2100 gnd vdd FILL
X_2231_ _2219_/Y _2227_/B gnd _2232_/A vdd NAND2X1
X_3280_ _3280_/A gnd _3280_/Y vdd INVX1
X_2300_ _2301_/A _2301_/B gnd _2300_/Y vdd NOR2X1
X_2093_ _2137_/Y gnd adrs_bus[7] vdd BUFX2
X_2162_ _2292_/B _2290_/B gnd _2167_/B vdd NAND2X1
XFILL71280x44100 gnd vdd FILL
X_2995_ gnd gnd _2995_/Y vdd INVX1
X_3616_ _3560_/B _3616_/B gnd _3617_/A vdd NAND2X1
X_3547_ _3559_/B gnd _3547_/Y vdd INVX1
X_4596_ _3550_/Y gnd _4596_/Y vdd INVX1
X_2429_ _2429_/A _2429_/B gnd _2429_/Y vdd XNOR2X1
X_3478_ _3513_/A _3513_/B _3477_/Y gnd _3481_/C vdd OAI21X1
X_4450_ _4450_/Q _4451_/CLK _4450_/D gnd vdd DFFPOSX1
X_2780_ _2776_/Y _2828_/A gnd _2788_/A vdd NOR2X1
X_4381_ _3816_/A _4383_/CLK _4381_/D gnd vdd DFFPOSX1
X_3401_ _3401_/A _3400_/Y _3401_/C gnd _3649_/B vdd NAND3X1
X_3332_ _3332_/A gnd _3334_/A vdd INVX1
X_3263_ _3263_/A _3341_/B _3262_/Y gnd _3263_/Y vdd OAI21X1
X_3194_ gnd _3194_/B _3194_/C gnd _3194_/Y vdd NAND3X1
X_2214_ _2195_/Y _2211_/Y _2214_/C gnd _2280_/A vdd OAI21X1
X_2145_ _2158_/A _4206_/A gnd _2145_/Y vdd NAND2X1
XSFILL14480x36100 gnd vdd FILL
X_2978_ _2978_/A _3346_/B _3346_/C gnd _2979_/A vdd NAND3X1
X_4579_ _4556_/C _4436_/CLK _4557_/Y gnd vdd DFFPOSX1
XSFILL29200x40100 gnd vdd FILL
X_3950_ _3950_/A _3950_/B _4027_/S gnd _3952_/A vdd MUX2X1
X_2763_ _2762_/A gnd _2765_/B vdd INVX1
X_2832_ _2832_/A _2101_/A _2766_/Y gnd _2836_/B vdd OAI21X1
X_2901_ _2901_/A _2900_/Y gnd _2901_/Y vdd NAND2X1
X_3881_ _3881_/A _3873_/B gnd _3882_/C vdd NOR2X1
X_4433_ _4433_/Q _4451_/CLK _4196_/Y gnd vdd DFFPOSX1
X_4502_ _4548_/C _4513_/B _4502_/C gnd _4504_/A vdd NAND3X1
X_2694_ _2690_/Y _2694_/B gnd _2703_/A vdd NAND2X1
X_4364_ _3714_/C _4300_/CLK _4364_/D gnd vdd DFFPOSX1
X_4295_ _3804_/A _4283_/B _4294_/Y gnd _4295_/Y vdd AOI21X1
X_3177_ gnd gnd _3178_/C vdd INVX1
X_3246_ gnd _3240_/B _3246_/C gnd _3248_/A vdd NAND3X1
X_3315_ _3313_/Y _3341_/B _3315_/C gnd _3315_/Y vdd OAI21X1
XSFILL29680x12100 gnd vdd FILL
X_2128_ _2140_/A _2126_/Y _2127_/Y gnd _2128_/Y vdd OAI21X1
X_4080_ _4343_/Q _4074_/S _4021_/C gnd _4081_/A vdd OAI21X1
X_3100_ _3098_/Y _3204_/B _3100_/C _3204_/D gnd _3100_/Y vdd OAI22X1
X_3031_ gnd _3343_/B gnd _3031_/Y vdd NAND2X1
X_3933_ _4314_/Q _4030_/S _3934_/C gnd _3934_/A vdd OAI21X1
X_2746_ _4072_/A _2660_/Y _2745_/Y _4050_/A gnd _2746_/Y vdd OAI22X1
X_3795_ _4208_/A _3802_/B gnd _3796_/C vdd NAND2X1
X_3864_ _4046_/A _3866_/B gnd _3865_/C vdd NAND2X1
X_2815_ _2488_/A gnd _2817_/A vdd INVX1
X_2677_ _2374_/A _2730_/A _2677_/C _4028_/A gnd _2678_/B vdd OAI22X1
X_4416_ _4416_/Q _4407_/CLK _4281_/Y gnd vdd DFFPOSX1
X_4347_ _4347_/Q _4345_/CLK _3780_/Y gnd vdd DFFPOSX1
XSFILL44720x10100 gnd vdd FILL
X_3229_ gnd gnd _3229_/Y vdd INVX1
X_4278_ _4415_/Q _4269_/B gnd _4278_/Y vdd NOR2X1
X_3580_ _4085_/A _3590_/B gnd _3582_/A vdd NAND2X1
X_2600_ _2600_/A _2600_/B gnd _2600_/Y vdd NAND2X1
X_4201_ _4418_/Q _3682_/A _4199_/B gnd _4204_/D vdd MUX2X1
X_2531_ _2351_/A _2530_/Y gnd _2533_/A vdd NAND2X1
X_2462_ _2606_/D gnd _2465_/A vdd INVX1
X_2393_ _2932_/B _4585_/B gnd _2396_/A vdd NOR2X1
X_4063_ _4241_/A _4390_/Q _4052_/S gnd _4063_/Y vdd MUX2X1
X_4132_ _3714_/C _4088_/B gnd _4132_/Y vdd NOR2X1
X_3014_ _3014_/A _3011_/Y _3014_/C gnd _3015_/B vdd NAND3X1
XSFILL14480x44100 gnd vdd FILL
X_3916_ _3649_/B gnd _3916_/Y vdd INVX1
X_3778_ _3811_/A _3802_/B _3777_/Y gnd _4346_/D vdd OAI21X1
X_3847_ _3813_/A _3846_/B _3847_/C gnd _3847_/Y vdd OAI21X1
X_2729_ _2721_/Y _2703_/Y _2728_/Y gnd _2729_/Y vdd AOI21X1
XBUFX2_insert161 _4435_/Q gnd _2252_/A vdd BUFX2
XBUFX2_insert194 _4454_/Q gnd _4072_/A vdd BUFX2
XBUFX2_insert172 _4432_/Q gnd _4184_/A vdd BUFX2
XBUFX2_insert183 _4429_/Q gnd _2890_/A vdd BUFX2
X_3563_ _3649_/A gnd _3563_/Y vdd INVX8
X_3632_ _3561_/B _3632_/CLK _3632_/D gnd vdd DFFPOSX1
XBUFX2_insert150 _4447_/Q gnd _2371_/A vdd BUFX2
X_3701_ _3771_/B _3700_/Y gnd _3704_/A vdd NOR2X1
X_2376_ _2374_/Y _2376_/B gnd _2385_/B vdd NOR2X1
X_2514_ _2514_/A _2514_/B gnd _3228_/A vdd AND2X2
X_4115_ _3877_/A _4124_/S _4111_/C gnd _4116_/A vdd OAI21X1
X_2445_ _2445_/A _2445_/B gnd _2445_/Y vdd XNOR2X1
X_3494_ _3494_/A _3508_/B _3508_/C gnd _3494_/Y vdd NAND3X1
X_4046_ _4046_/A _3932_/B gnd _4046_/Y vdd NOR2X1
XSFILL45040x8100 gnd vdd FILL
X_2230_ _2229_/Y gnd _2230_/Y vdd INVX1
X_2161_ _2151_/A _2159_/Y _2160_/Y gnd _2161_/Y vdd OAI21X1
X_2092_ _2092_/A gnd adrs_bus[6] vdd BUFX2
X_2994_ _2441_/Y gnd _2994_/Y vdd INVX1
X_3615_ _3614_/Y _3573_/B _3615_/C gnd _3630_/D vdd AOI21X1
X_4595_ _4594_/A _4593_/Y _4594_/Y gnd _4595_/Y vdd OAI21X1
X_3546_ _4628_/A _3546_/B gnd _3546_/Y vdd NOR2X1
X_2428_ _2428_/A _2127_/B gnd _2428_/Y vdd XNOR2X1
X_3477_ _3172_/Y gnd _3477_/Y vdd INVX1
X_2359_ _2428_/A _2127_/B gnd _3089_/A vdd AND2X2
X_4029_ _4027_/Y _4207_/B _4028_/Y gnd _4450_/D vdd AOI21X1
XSFILL29200x38100 gnd vdd FILL
X_3331_ _3331_/A _2950_/B _3331_/C _3201_/D gnd _3335_/B vdd OAI22X1
X_4380_ _3814_/A _4383_/CLK _4380_/D gnd vdd DFFPOSX1
X_3400_ _2965_/B _3410_/A _3400_/C gnd _3400_/Y vdd OAI21X1
X_2144_ _4575_/Q gnd _2144_/Y vdd INVX1
X_3193_ _3193_/A _3141_/B gnd _3196_/B vdd NAND2X1
X_3262_ gnd _3340_/B gnd _3262_/Y vdd NAND2X1
X_2213_ _2209_/Y _2213_/B _2207_/Y gnd _2214_/C vdd AOI21X1
XFILL71120x2100 gnd vdd FILL
XSFILL14480x52100 gnd vdd FILL
X_2977_ _2290_/Y _2977_/B _3194_/B gnd _2977_/Y vdd NAND3X1
X_4578_ _4578_/Q _4436_/CLK _4551_/Y gnd vdd DFFPOSX1
X_3529_ _3528_/Y _3508_/B _3508_/C gnd _3529_/Y vdd NAND3X1
XFILL71280x8100 gnd vdd FILL
XSFILL14640x12100 gnd vdd FILL
XSFILL44560x48100 gnd vdd FILL
X_2900_ _2898_/Y _2895_/A _2896_/A _2900_/D gnd _2900_/Y vdd AOI22X1
X_2762_ _2762_/A _2762_/B _2762_/C _2762_/D gnd _2766_/A vdd OAI22X1
X_2831_ _2831_/A _2831_/B _2831_/C gnd _2837_/A vdd OAI21X1
X_3880_ _3813_/A _3896_/B _3879_/Y gnd _4331_/D vdd AOI21X1
X_4501_ _4495_/A _4501_/B _4495_/B gnd _4513_/B vdd NAND3X1
X_4294_ _4423_/Q _4283_/B gnd _4294_/Y vdd NOR2X1
X_4432_ _4432_/Q _4451_/CLK _4432_/D gnd vdd DFFPOSX1
XSFILL44240x30100 gnd vdd FILL
X_4363_ _4363_/Q _4345_/CLK _3713_/Y gnd vdd DFFPOSX1
X_3314_ gnd _3340_/B gnd _3315_/C vdd NAND2X1
X_2693_ _2724_/B _2693_/B _2693_/C _2881_/D gnd _2694_/B vdd AOI22X1
X_3176_ _3176_/A gnd _3178_/A vdd INVX1
X_2127_ _2140_/A _2127_/B gnd _2127_/Y vdd NAND2X1
X_3245_ _3245_/A _3141_/B gnd _3248_/B vdd NAND2X1
X_3030_ _3030_/A _3029_/Y gnd _3042_/B vdd NOR2X1
X_3863_ _3729_/A _3862_/B _3863_/C gnd _3863_/Y vdd OAI21X1
X_3932_ _3932_/A _3932_/B gnd _3932_/Y vdd NOR2X1
X_3794_ _3794_/A _3803_/B _3793_/Y gnd _3794_/Y vdd OAI21X1
X_2676_ _2676_/A gnd _2677_/C vdd INVX1
X_2745_ _2745_/A gnd _2745_/Y vdd INVX1
X_2814_ _2810_/Y _2813_/Y gnd _2814_/Y vdd NOR2X1
X_4346_ _4109_/A _4345_/CLK _4346_/D gnd vdd DFFPOSX1
X_4415_ _4415_/Q _4394_/CLK _4279_/Y gnd vdd DFFPOSX1
X_4277_ _3752_/A _4277_/B _4276_/Y gnd _4414_/D vdd AOI21X1
X_3228_ _3228_/A gnd _3230_/A vdd INVX1
X_3159_ _3159_/A _3341_/B _3159_/C gnd _3160_/B vdd OAI21X1
XSFILL29520x100 gnd vdd FILL
XSFILL29200x46100 gnd vdd FILL
X_2530_ _2351_/B gnd _2530_/Y vdd INVX1
X_4200_ _4200_/A _4198_/Y _4199_/C _4200_/D gnd _4205_/B vdd OAI22X1
X_2461_ _2474_/D _2461_/B gnd _2461_/Y vdd XNOR2X1
X_4131_ _4131_/A _3814_/A _4153_/S gnd _4131_/Y vdd MUX2X1
X_2392_ _2932_/B _2392_/B gnd _2392_/Y vdd AND2X2
X_4062_ _4062_/A _4040_/B _4061_/Y gnd _4453_/D vdd AOI21X1
X_3013_ _3143_/A gnd gnd _3143_/D gnd _3014_/C vdd AOI22X1
X_3846_ _3947_/A _3846_/B gnd _3847_/C vdd NAND2X1
X_3915_ _3914_/Y _3915_/B _4027_/S gnd _3919_/A vdd MUX2X1
X_2659_ _2659_/A _2659_/B gnd _2659_/Y vdd NAND2X1
X_3777_ _4109_/A _3802_/B gnd _3777_/Y vdd NAND2X1
X_2728_ _2723_/Y _2703_/A _2727_/Y gnd _2728_/Y vdd OAI21X1
XSFILL29680x18100 gnd vdd FILL
X_4329_ _4329_/Q _4394_/CLK _3876_/Y gnd vdd DFFPOSX1
XSFILL14640x20100 gnd vdd FILL
XBUFX2_insert140 _3917_/Y gnd _4207_/B vdd BUFX2
XBUFX2_insert151 _4438_/Q gnd _2762_/C vdd BUFX2
X_3700_ _3771_/A gnd _3700_/Y vdd INVX1
XBUFX2_insert162 _4435_/Q gnd _2374_/B vdd BUFX2
XBUFX2_insert173 _4432_/Q gnd _2782_/A vdd BUFX2
XBUFX2_insert195 _4454_/Q gnd _2102_/A vdd BUFX2
X_2513_ _2510_/Y _2511_/Y gnd _2514_/A vdd OR2X2
X_3631_ _3560_/B _4431_/CLK _3631_/D gnd vdd DFFPOSX1
XBUFX2_insert184 _4429_/Q gnd _2190_/A vdd BUFX2
X_3493_ data_in[9] gnd _3494_/A vdd INVX1
X_3562_ _3562_/A _3553_/A gnd _4626_/A vdd AND2X2
X_2375_ _4028_/A _4206_/A gnd _2376_/B vdd XOR2X1
X_4114_ _3936_/A _4180_/B gnd _4116_/B vdd NOR2X1
X_2444_ _2614_/C _2104_/A gnd _2445_/B vdd XNOR2X1
X_4045_ _4045_/A _3688_/A _4036_/B gnd _4045_/Y vdd MUX2X1
XSFILL44720x16100 gnd vdd FILL
X_3829_ _3729_/A _3823_/B _3828_/Y gnd _3829_/Y vdd AOI21X1
X_2160_ _2151_/A _4261_/A gnd _2160_/Y vdd NAND2X1
XSFILL59760x32100 gnd vdd FILL
X_2091_ _2091_/A gnd adrs_bus[5] vdd BUFX2
X_3614_ _3559_/B _3605_/B gnd _3614_/Y vdd NAND2X1
X_2993_ _2991_/Y _2950_/B _2992_/Y _3201_/D gnd _2997_/B vdd OAI22X1
X_2427_ _2427_/A _2427_/B _2427_/C _2427_/D gnd _2430_/C vdd AOI22X1
X_3476_ _3422_/B _4602_/A gnd _3476_/Y vdd NAND2X1
X_4594_ _4594_/A _2127_/B gnd _4594_/Y vdd NAND2X1
X_3545_ _3545_/A gnd _3546_/B vdd INVX1
X_4028_ _4028_/A _4207_/B _4206_/C gnd _4028_/Y vdd OAI21X1
X_2289_ _2289_/A _2289_/B gnd _3371_/A vdd NAND2X1
X_2358_ _2301_/A _2301_/B gnd _2358_/Y vdd AND2X2
XSFILL59440x4100 gnd vdd FILL
XSFILL14160x32100 gnd vdd FILL
X_3330_ gnd gnd _3331_/C vdd INVX1
X_2143_ _2158_/A _2141_/Y _2143_/C gnd _2143_/Y vdd OAI21X1
X_3192_ _3187_/Y _3192_/B _3191_/Y gnd _3197_/A vdd NAND3X1
X_3261_ gnd gnd _3263_/A vdd INVX1
XSFILL44240x28100 gnd vdd FILL
X_2212_ _2199_/Y _2211_/Y gnd _2215_/A vdd NOR2X1
X_4577_ _2150_/A _4451_/CLK _4544_/Y gnd vdd DFFPOSX1
XSFILL29680x26100 gnd vdd FILL
X_2976_ _2293_/Y _3090_/B _3110_/C gnd _2976_/Y vdd NAND3X1
X_3528_ data_in[14] gnd _3528_/Y vdd INVX1
X_3459_ _3458_/Y _3508_/B _3508_/C gnd _3459_/Y vdd NAND3X1
XSFILL59280x44100 gnd vdd FILL
XSFILL29360x8100 gnd vdd FILL
X_2830_ _2830_/A _2830_/B _2784_/Y gnd _2831_/A vdd OAI21X1
XSFILL44560x2100 gnd vdd FILL
X_2761_ _2761_/A gnd _2762_/D vdd INVX1
X_4500_ _4493_/C _4489_/C _4499_/Y gnd _4502_/C vdd OAI21X1
X_2692_ _2880_/A gnd _2693_/C vdd INVX1
X_4431_ _4431_/Q _4431_/CLK _4431_/D gnd vdd DFFPOSX1
X_3244_ _3244_/A _3240_/Y _3244_/C gnd _3249_/A vdd NAND3X1
X_4293_ _3902_/A _4292_/B _4293_/C gnd _4293_/Y vdd AOI21X1
X_4362_ _3932_/A _4345_/CLK _3711_/Y gnd vdd DFFPOSX1
X_3313_ gnd gnd _3313_/Y vdd INVX1
X_3175_ _3175_/A _2950_/B _3175_/C _3201_/D gnd _3179_/B vdd OAI22X1
X_2126_ _4488_/B gnd _2126_/Y vdd INVX1
X_2959_ gnd gnd _2959_/Y vdd INVX1
XSFILL44720x24100 gnd vdd FILL
XSFILL59760x40100 gnd vdd FILL
X_3862_ _3862_/A _3862_/B gnd _3863_/C vdd NAND2X1
X_3931_ _4109_/A _4378_/Q _4030_/S gnd _3934_/D vdd MUX2X1
X_2813_ _2881_/B _2813_/B _2813_/C _2881_/D gnd _2813_/Y vdd OAI22X1
X_3793_ _4354_/Q _3803_/B gnd _3793_/Y vdd NAND2X1
X_2675_ _2374_/B gnd _2730_/A vdd INVX1
X_2744_ _2744_/A _2729_/Y _2744_/C gnd _2759_/B vdd OAI21X1
XSFILL14480x6100 gnd vdd FILL
X_4414_ _4276_/A _4394_/CLK _4414_/D gnd vdd DFFPOSX1
X_3227_ _3227_/A _2950_/B _3226_/Y _3201_/D gnd _3231_/B vdd OAI22X1
X_4345_ _4345_/Q _4345_/CLK _3776_/Y gnd vdd DFFPOSX1
XFILL71120x8100 gnd vdd FILL
X_4276_ _4276_/A _4277_/B gnd _4276_/Y vdd NOR2X1
X_3158_ gnd _3340_/B gnd _3159_/C vdd NAND2X1
X_2109_ _2881_/B gnd data_out[7] vdd BUFX2
X_3089_ _3089_/A _3141_/B gnd _3092_/B vdd NAND2X1
XSFILL14160x40100 gnd vdd FILL
XBUFX2_insert300 _4425_/Q gnd _2392_/B vdd BUFX2
XSFILL14640x18100 gnd vdd FILL
X_2460_ _2606_/D _2465_/B gnd _2461_/B vdd XOR2X1
X_4061_ _4061_/A _4040_/B _4239_/C gnd _4061_/Y vdd OAI21X1
X_2391_ _2391_/A _2390_/Y gnd _2391_/Y vdd NOR2X1
X_4130_ _4130_/A _4130_/B _4129_/Y gnd _4427_/D vdd AOI21X1
X_3012_ gnd _3240_/B _3246_/C gnd _3014_/A vdd NAND3X1
X_3845_ _3811_/A _3866_/B _3845_/C gnd _4298_/D vdd OAI21X1
X_3776_ _3843_/A _3775_/B _3776_/C gnd _3776_/Y vdd OAI21X1
X_3914_ _3913_/Y _3914_/B _3982_/C _3914_/D gnd _3914_/Y vdd OAI22X1
X_2589_ _2588_/Y _2786_/A _2786_/C _2586_/Y gnd _2642_/C vdd AOI22X1
X_2658_ _2569_/A gnd _2659_/B vdd INVX1
XSFILL29680x34100 gnd vdd FILL
X_2727_ _2726_/Y _2727_/B _2727_/C gnd _2727_/Y vdd AOI21X1
X_4259_ _4259_/A _4257_/Y _4199_/C _4259_/D gnd _4260_/A vdd OAI22X1
X_4328_ _3873_/A _4297_/CLK _4328_/D gnd vdd DFFPOSX1
XSFILL59280x52100 gnd vdd FILL
XBUFX2_insert141 _3917_/Y gnd _4240_/B vdd BUFX2
XBUFX2_insert174 _4432_/Q gnd _2875_/A vdd BUFX2
XBUFX2_insert152 _4438_/Q gnd _2571_/B vdd BUFX2
XBUFX2_insert163 _4263_/Y gnd _4269_/B vdd BUFX2
XBUFX2_insert185 _4429_/Q gnd _2488_/A vdd BUFX2
X_3630_ _3559_/B _3632_/CLK _3630_/D gnd vdd DFFPOSX1
XBUFX2_insert130 _3410_/Y gnd _3434_/A vdd BUFX2
X_2512_ _2511_/Y _2510_/Y gnd _2514_/B vdd NAND2X1
X_3492_ _3513_/A _3513_/B _3492_/C gnd _3492_/Y vdd OAI21X1
X_2443_ _2443_/A _2443_/B _2442_/Y gnd _2445_/A vdd AOI21X1
XBUFX2_insert196 _3409_/Y gnd _2124_/A vdd BUFX2
X_3561_ _3561_/A _3561_/B gnd _4623_/A vdd AND2X2
X_2374_ _2374_/A _2374_/B gnd _2374_/Y vdd XOR2X1
X_4044_ _4043_/Y _4044_/B _4004_/C _4041_/Y gnd _4049_/B vdd OAI22X1
X_4113_ _3935_/A _3935_/B _4124_/S gnd _4113_/Y vdd MUX2X1
X_3759_ _4199_/A _3760_/B gnd _3759_/Y vdd NAND2X1
X_3828_ _4208_/B _3823_/B gnd _3828_/Y vdd NOR2X1
XSFILL44720x32100 gnd vdd FILL
X_2090_ _2128_/Y gnd adrs_bus[4] vdd BUFX2
X_2992_ gnd gnd _2992_/Y vdd INVX1
X_3613_ _3612_/Y _3613_/B _3570_/C gnd _3629_/D vdd AOI21X1
X_4593_ _4593_/A gnd _4593_/Y vdd INVX1
X_2426_ _2382_/A _4195_/A gnd _2427_/D vdd OR2X2
X_3475_ _3469_/Y _3474_/Y gnd _3475_/Y vdd NAND2X1
X_3544_ _3561_/A _3544_/B gnd _3441_/B vdd NOR2X1
X_4027_ _4026_/Y _4027_/B _4027_/S gnd _4027_/Y vdd MUX2X1
X_2288_ _2288_/A _2288_/B gnd _2289_/B vdd NAND2X1
X_2357_ _2298_/A _2298_/B gnd _2357_/Y vdd AND2X2
X_3260_ _3260_/A _3130_/B _3260_/C _3130_/D gnd _3264_/A vdd OAI22X1
X_2142_ _2158_/A _4195_/A gnd _2143_/C vdd NAND2X1
X_3191_ _3190_/Y _3191_/B gnd _3191_/Y vdd AND2X2
X_2211_ _2206_/B _2209_/Y gnd _2211_/Y vdd NAND2X1
XSFILL44240x44100 gnd vdd FILL
X_2975_ _2986_/A _2986_/B gnd _2975_/Y vdd NOR2X1
X_4576_ _2147_/A _4436_/CLK _4576_/D gnd vdd DFFPOSX1
X_3527_ _3513_/A _3513_/B _3527_/C gnd _3527_/Y vdd OAI21X1
XSFILL29680x42100 gnd vdd FILL
X_2409_ _4072_/A _4250_/A gnd _2415_/B vdd XNOR2X1
X_3458_ data_in[4] gnd _3458_/Y vdd INVX1
X_3389_ _2986_/A _3382_/Y gnd _3389_/Y vdd NAND2X1
XSFILL60240x26100 gnd vdd FILL
X_2760_ _2849_/A gnd _2762_/B vdd INVX1
X_2691_ _2881_/B gnd _2724_/B vdd INVX1
X_4430_ _4430_/Q _4431_/CLK _4430_/D gnd vdd DFFPOSX1
X_4292_ _4292_/A _4292_/B gnd _4293_/C vdd NOR2X1
X_3243_ _3242_/Y _3243_/B gnd _3244_/C vdd AND2X2
X_3312_ _3310_/Y _3130_/B _3312_/C _3130_/D gnd _3312_/Y vdd OAI22X1
X_4361_ _3921_/A _4345_/CLK _3709_/Y gnd vdd DFFPOSX1
X_3174_ gnd gnd _3175_/C vdd INVX1
X_2125_ _2124_/A _2123_/Y _2125_/C gnd _2089_/A vdd OAI21X1
XSFILL59440x20100 gnd vdd FILL
X_2958_ gnd gnd _2963_/A vdd INVX1
X_4559_ _2159_/A gnd _4559_/Y vdd INVX1
X_4628_ _4628_/A _4626_/Y _4627_/Y gnd _4628_/Y vdd OAI21X1
X_2889_ _2190_/B gnd _2889_/Y vdd INVX1
XSFILL14160x38100 gnd vdd FILL
X_3930_ _3930_/A _3951_/B _3929_/Y gnd _4441_/D vdd AOI21X1
X_3861_ _3794_/A _3870_/B _3860_/Y gnd _4306_/D vdd OAI21X1
X_2743_ _2671_/Y _2743_/B _2743_/C gnd _2744_/C vdd AOI21X1
X_3792_ _4283_/A _3792_/B _3791_/Y gnd _4353_/D vdd OAI21X1
X_2812_ _2880_/A gnd _2813_/C vdd INVX1
X_2674_ _2374_/B _2731_/B _2676_/A _2674_/D gnd _2734_/C vdd OAI22X1
X_4413_ _4274_/A _4383_/CLK _4413_/D gnd vdd DFFPOSX1
X_4344_ _3773_/A _4345_/CLK _4344_/D gnd vdd DFFPOSX1
X_3226_ gnd gnd _3226_/Y vdd INVX1
X_3157_ gnd gnd _3159_/A vdd INVX1
X_4275_ _3717_/A _4277_/B _4274_/Y gnd _4413_/D vdd AOI21X1
X_2108_ _2881_/D gnd data_out[6] vdd BUFX2
XSFILL29200x8100 gnd vdd FILL
X_3088_ _3088_/A _3084_/Y _3087_/Y gnd _3088_/Y vdd NAND3X1
XSFILL44400x2100 gnd vdd FILL
XSFILL14640x34100 gnd vdd FILL
XBUFX2_insert301 _4425_/Q gnd _2752_/A vdd BUFX2
XSFILL44080x2100 gnd vdd FILL
X_4060_ _4060_/A _4055_/Y _4027_/S gnd _4062_/A vdd MUX2X1
X_2390_ _2428_/A _2892_/A gnd _2390_/Y vdd XOR2X1
X_3011_ _2356_/Y _3141_/B gnd _3011_/Y vdd NAND2X1
X_3913_ _3873_/A _3992_/B _3982_/C gnd _3913_/Y vdd OAI21X1
XSFILL44240x52100 gnd vdd FILL
X_3844_ _3936_/A _3866_/B gnd _3845_/C vdd NAND2X1
X_3775_ _4345_/Q _3775_/B gnd _3776_/C vdd NAND2X1
X_2726_ _2880_/A _2690_/D gnd _2726_/Y vdd NOR2X1
X_4327_ _4327_/Q _4359_/CLK _3770_/Y gnd vdd DFFPOSX1
X_2588_ _2318_/B gnd _2588_/Y vdd INVX1
X_2657_ _2569_/A _2758_/B gnd _2657_/Y vdd NAND2X1
XSFILL29680x50100 gnd vdd FILL
X_4258_ _4343_/Q _4252_/S _4199_/C gnd _4259_/A vdd OAI21X1
X_4189_ _4189_/A _4187_/Y _4254_/C _4186_/Y gnd _4189_/Y vdd OAI22X1
X_3209_ gnd gnd _3211_/A vdd INVX1
XSFILL14320x6100 gnd vdd FILL
XSFILL59760x46100 gnd vdd FILL
XBUFX2_insert142 _3917_/Y gnd _4040_/B vdd BUFX2
XBUFX2_insert120 _3642_/Q gnd _4199_/C vdd BUFX2
XBUFX2_insert197 _3409_/Y gnd _2158_/A vdd BUFX2
XBUFX2_insert153 _4438_/Q gnd _4250_/A vdd BUFX2
XBUFX2_insert175 _4432_/Q gnd _2421_/B vdd BUFX2
XBUFX2_insert164 _4263_/Y gnd _4287_/B vdd BUFX2
X_3560_ _4628_/A _3560_/B gnd _4620_/A vdd AND2X2
XBUFX2_insert131 _3421_/Q gnd _3601_/A vdd BUFX2
XBUFX2_insert186 _4429_/Q gnd _4597_/B vdd BUFX2
X_2511_ _2778_/A _2098_/A gnd _2511_/Y vdd XNOR2X1
X_3491_ _3491_/A gnd _3492_/C vdd INVX1
X_2442_ _2442_/A _2442_/B gnd _2442_/Y vdd NOR2X1
X_2373_ _2371_/Y _2372_/Y gnd _2373_/Y vdd NOR2X1
X_4043_ _4221_/A _4036_/B _4004_/C gnd _4043_/Y vdd OAI21X1
X_4112_ _4112_/A _4112_/B _4111_/C _4112_/D gnd _4117_/B vdd OAI22X1
X_3827_ _3794_/A _3832_/B _3826_/Y gnd _4386_/D vdd AOI21X1
X_3758_ _4283_/A _3760_/B _3758_/C gnd _4321_/D vdd OAI21X1
X_3689_ _3764_/A _3685_/B _3689_/C gnd _4404_/D vdd AOI21X1
X_2709_ _2717_/B _2609_/A _2708_/Y _2899_/A gnd _2756_/B vdd AOI22X1
XSFILL14160x46100 gnd vdd FILL
X_2991_ _2991_/A gnd _2991_/Y vdd INVX1
X_3612_ _3545_/A _3616_/B gnd _3612_/Y vdd NAND2X1
X_3543_ _3557_/B gnd _3544_/B vdd INVX1
X_4592_ _4594_/A _4592_/B _4591_/Y gnd _4592_/Y vdd OAI21X1
X_2425_ _2382_/A _2682_/A gnd _2427_/C vdd NAND2X1
X_3474_ _3495_/A _3473_/Y _3474_/C gnd _3474_/Y vdd NAND3X1
X_2356_ _2295_/A _2295_/B gnd _2356_/Y vdd AND2X2
X_4026_ _4025_/Y _4024_/Y _4010_/C _4026_/D gnd _4026_/Y vdd OAI22X1
X_2287_ _2287_/A _2287_/B _2272_/B gnd _2288_/B vdd OAI21X1
XSFILL29360x22100 gnd vdd FILL
XSFILL14640x42100 gnd vdd FILL
X_3190_ gnd _3346_/B _3346_/C gnd _3190_/Y vdd NAND3X1
X_2210_ _2206_/Y _2209_/Y gnd _2210_/Y vdd XNOR2X1
X_2141_ _4574_/Q gnd _2141_/Y vdd INVX1
XSFILL59440x18100 gnd vdd FILL
X_2974_ gnd _3343_/B gnd _2980_/A vdd NAND2X1
X_4575_ _4575_/Q _4436_/CLK _4531_/Y gnd vdd DFFPOSX1
X_3526_ _3526_/A gnd _3527_/C vdd INVX1
XSFILL44720x38100 gnd vdd FILL
X_2408_ _2848_/A _4261_/A gnd _2415_/A vdd XNOR2X1
X_3388_ _3388_/A gnd _3390_/B vdd INVX1
X_3457_ _3513_/A _3513_/B _3456_/Y gnd _3460_/C vdd OAI21X1
X_2339_ _2429_/A _2433_/A gnd _2339_/Y vdd OR2X2
X_4009_ _4187_/A _4020_/B gnd _4011_/B vdd NOR2X1
XSFILL44400x20100 gnd vdd FILL
XFILL71120x22100 gnd vdd FILL
X_3311_ gnd gnd _3312_/C vdd INVX1
X_2690_ _2690_/A _2881_/B _2880_/A _2690_/D gnd _2690_/Y vdd AOI22X1
X_4360_ _4360_/Q _4345_/CLK _3707_/Y gnd vdd DFFPOSX1
X_4291_ _3692_/A _4292_/B _4290_/Y gnd _4291_/Y vdd AOI21X1
X_3173_ _3173_/A gnd _3175_/A vdd INVX1
X_3242_ gnd _3294_/B _3268_/C gnd _3242_/Y vdd NAND3X1
X_2124_ _2124_/A _4591_/B gnd _2125_/C vdd NAND2X1
X_4627_ _4628_/A _4261_/A gnd _4627_/Y vdd NAND2X1
X_2957_ _2957_/A _2950_/Y gnd _2957_/Y vdd NOR2X1
X_2888_ _2914_/A _2190_/B _2428_/A _2887_/Y gnd _2893_/C vdd AOI22X1
X_4558_ _4628_/Y _4558_/B gnd _4558_/Y vdd NAND2X1
X_4489_ _4548_/C _4486_/Y _4489_/C gnd _4489_/Y vdd NAND3X1
X_3509_ _3495_/A _3508_/Y _3509_/C gnd _3509_/Y vdd NAND3X1
X_3860_ _4024_/A _3870_/B gnd _3860_/Y vdd NAND2X1
X_2742_ _2742_/A _2740_/Y _2748_/A gnd _2743_/C vdd OAI21X1
X_3791_ _4186_/A _3792_/B gnd _3791_/Y vdd NAND2X1
X_2811_ _2693_/B gnd _2813_/B vdd INVX1
XSFILL14320x14100 gnd vdd FILL
X_2673_ _2673_/A gnd _2674_/D vdd INVX1
X_4343_ _4343_/Q _4359_/CLK _3904_/Y gnd vdd DFFPOSX1
X_4274_ _4274_/A _4277_/B gnd _4274_/Y vdd NOR2X1
X_4412_ _4412_/Q _4394_/CLK _4412_/D gnd vdd DFFPOSX1
X_3225_ _3225_/A gnd _3227_/A vdd INVX1
X_3156_ _3156_/A _3130_/B _3155_/Y _3130_/D gnd _3160_/A vdd OAI22X1
X_2107_ _2723_/B gnd data_out[5] vdd BUFX2
X_3087_ _3087_/A _3085_/Y gnd _3087_/Y vdd AND2X2
XSFILL29680x48100 gnd vdd FILL
X_3989_ _3989_/A _3989_/B _3988_/C _3989_/D gnd _3994_/B vdd OAI22X1
XSFILL29360x30100 gnd vdd FILL
XSFILL14640x50100 gnd vdd FILL
X_3010_ _3005_/Y _3006_/Y _3010_/C gnd _3015_/A vdd NAND3X1
X_3843_ _3843_/A _3846_/B _3842_/Y gnd _4297_/D vdd OAI21X1
X_3912_ _3840_/A _3943_/B gnd _3914_/B vdd NOR2X1
X_2656_ _2659_/A gnd _2758_/B vdd INVX1
X_2725_ _2693_/B _2724_/B gnd _2727_/B vdd NAND2X1
X_3774_ _3740_/A _3775_/B _3773_/Y gnd _4344_/D vdd OAI21X1
X_4257_ _3870_/A _4198_/B gnd _4257_/Y vdd NOR2X1
X_2587_ _2586_/Y _2786_/C gnd _2590_/C vdd OR2X2
X_4326_ _3767_/A _4407_/CLK _4326_/D gnd vdd DFFPOSX1
XSFILL14800x10100 gnd vdd FILL
X_4188_ _4010_/A _4199_/B _4254_/C gnd _4189_/A vdd OAI21X1
X_3208_ _3208_/A _3130_/B _3208_/C _3130_/D gnd _3212_/A vdd OAI22X1
X_3139_ _3139_/A _3137_/Y gnd _3139_/Y vdd AND2X2
XBUFX2_insert110 _4452_/Q gnd _4050_/A vdd BUFX2
XBUFX2_insert154 _4438_/Q gnd _2572_/A vdd BUFX2
X_2510_ _2509_/Y _2500_/B _2508_/Y gnd _2510_/Y vdd OAI21X1
XBUFX2_insert121 _3642_/Q gnd _4247_/C vdd BUFX2
XBUFX2_insert198 _3409_/Y gnd _2140_/A vdd BUFX2
X_3490_ _3532_/A _3490_/B gnd _3496_/A vdd NAND2X1
XBUFX2_insert143 _3649_/Y gnd _3703_/B vdd BUFX2
XSFILL58960x4100 gnd vdd FILL
XBUFX2_insert132 _3421_/Q gnd _3575_/A vdd BUFX2
XBUFX2_insert187 _4429_/Q gnd _2394_/B vdd BUFX2
XBUFX2_insert176 _3625_/Q gnd _3561_/A vdd BUFX2
XBUFX2_insert165 _4263_/Y gnd _4277_/B vdd BUFX2
X_4111_ _4314_/Q _4124_/S _4111_/C gnd _4112_/A vdd OAI21X1
X_2441_ _2441_/A _2443_/A gnd _2441_/Y vdd XNOR2X1
XSFILL15120x2100 gnd vdd FILL
X_2372_ _2418_/A _4600_/B gnd _2372_/Y vdd XOR2X1
X_4042_ _4042_/A _3932_/B gnd _4044_/B vdd NOR2X1
X_3826_ _3826_/A _3832_/B gnd _3826_/Y vdd NOR2X1
X_2639_ _2779_/B gnd _2640_/A vdd INVX1
X_3757_ _4010_/A _3760_/B gnd _3758_/C vdd NAND2X1
X_3688_ _3688_/A _3685_/B gnd _3689_/C vdd NOR2X1
X_2708_ _2896_/A gnd _2708_/Y vdd INVX1
X_4309_ _4057_/A _4298_/CLK _4309_/D gnd vdd DFFPOSX1
XSFILL59920x22100 gnd vdd FILL
X_2990_ _2957_/Y _2990_/B _2990_/C gnd _3424_/A vdd NAND3X1
X_3611_ _3610_/Y _3611_/B _3579_/C gnd _3611_/Y vdd AOI21X1
X_3473_ _3472_/Y _3508_/B _3508_/C gnd _3473_/Y vdd NAND3X1
X_3542_ _3562_/A _3541_/Y gnd _4584_/A vdd NOR2X1
X_4591_ _4594_/A _4591_/B gnd _4591_/Y vdd NAND2X1
X_2286_ _2272_/Y gnd _2287_/A vdd INVX1
X_2424_ _4061_/A _2665_/A gnd _2427_/A vdd OR2X2
X_2355_ _2429_/A _2433_/A gnd _2355_/Y vdd AND2X2
X_4025_ _4025_/A _4012_/S _4010_/C gnd _4025_/Y vdd OAI21X1
X_3809_ _3843_/A _3809_/B _3808_/Y gnd _3809_/Y vdd AOI21X1
XSFILL44400x18100 gnd vdd FILL
XSFILL29840x16100 gnd vdd FILL
X_2140_ _2140_/A _2138_/Y _2139_/Y gnd _2140_/Y vdd OAI21X1
XSFILL43760x46100 gnd vdd FILL
X_2973_ _3372_/C _2977_/B gnd _3343_/B vdd AND2X2
XSFILL59440x34100 gnd vdd FILL
X_4574_ _4574_/Q _4436_/CLK _4574_/D gnd vdd DFFPOSX1
X_3525_ _3518_/A _4623_/A gnd _3531_/A vdd NAND2X1
X_3456_ _3094_/Y gnd _3456_/Y vdd INVX1
X_4008_ _4186_/A _4186_/B _4012_/S gnd _4008_/Y vdd MUX2X1
X_2269_ _2255_/Y _2264_/Y _2268_/Y gnd _2287_/B vdd AOI21X1
X_2338_ _2336_/Y _2337_/Y gnd _3370_/A vdd NOR2X1
X_3387_ _3410_/B _3387_/B _3416_/A gnd _2112_/A vdd OAI21X1
X_2407_ _2407_/A _2406_/Y gnd _2407_/Y vdd NAND2X1
X_4290_ _4056_/A _4292_/B gnd _4290_/Y vdd NOR2X1
X_3310_ gnd gnd _3310_/Y vdd INVX1
X_3241_ _3241_/A _2961_/A _3267_/C gnd _3243_/B vdd NAND3X1
X_3172_ _3153_/Y _3172_/B _3171_/Y gnd _3172_/Y vdd NAND3X1
X_2123_ _4488_/A gnd _2123_/Y vdd INVX1
X_2956_ _2951_/Y _3204_/B _2956_/C _3204_/D gnd _2957_/A vdd OAI22X1
X_2887_ _2892_/A gnd _2887_/Y vdd INVX1
X_4626_ _4626_/A gnd _4626_/Y vdd INVX1
X_4557_ _4555_/Y _4556_/Y _4557_/C gnd _4557_/Y vdd AOI21X1
X_4488_ _4488_/A _4488_/B _4488_/C gnd _4489_/C vdd NAND3X1
X_3508_ _3507_/Y _3508_/B _3508_/C gnd _3508_/Y vdd NAND3X1
X_3439_ _3495_/A _3438_/Y _3436_/Y gnd _3439_/Y vdd NAND3X1
XSFILL59920x30100 gnd vdd FILL
XSFILL29360x28100 gnd vdd FILL
XFILL70960x44100 gnd vdd FILL
XSFILL14640x48100 gnd vdd FILL
X_2672_ _2829_/B gnd _2731_/B vdd INVX1
X_2741_ _2660_/Y _4072_/A _2670_/A gnd _2742_/A vdd OAI21X1
X_3790_ _4281_/A _3792_/B _3789_/Y gnd _3790_/Y vdd OAI21X1
X_4411_ _4124_/A _4298_/CLK _4411_/D gnd vdd DFFPOSX1
X_2810_ _2482_/A _2822_/B _2916_/A _2810_/D gnd _2810_/Y vdd OAI22X1
X_4342_ _4069_/A _4417_/CLK _4342_/D gnd vdd DFFPOSX1
X_3224_ _3224_/A _3212_/Y _3223_/Y gnd _3491_/A vdd NAND3X1
XSFILL14320x30100 gnd vdd FILL
X_4273_ _4273_/A _4269_/B _4273_/C gnd _4412_/D vdd AOI21X1
.ends

