magic
tech scmos
magscale 1 2
timestamp 1596033377
<< metal1 >>
rect 2938 5414 2950 5416
rect 5946 5414 5958 5416
rect 2923 5406 2925 5414
rect 2933 5406 2935 5414
rect 2943 5406 2945 5414
rect 2953 5406 2955 5414
rect 2963 5406 2965 5414
rect 5931 5406 5933 5414
rect 5941 5406 5943 5414
rect 5951 5406 5953 5414
rect 5961 5406 5963 5414
rect 5971 5406 5973 5414
rect 2938 5404 2950 5406
rect 5946 5404 5958 5406
rect 2280 5376 2284 5384
rect 829 5357 844 5363
rect 269 5337 284 5343
rect 365 5337 380 5343
rect 877 5343 883 5363
rect 1117 5357 1139 5363
rect 3373 5357 3395 5363
rect 3501 5357 3523 5363
rect 3933 5357 3971 5363
rect 4605 5357 4643 5363
rect 6205 5357 6243 5363
rect 7005 5357 7043 5363
rect 804 5337 835 5343
rect 877 5337 908 5343
rect 1581 5337 1596 5343
rect 2477 5337 2499 5343
rect 3956 5337 3987 5343
rect 5037 5337 5052 5343
rect 5436 5343 5444 5348
rect 5421 5337 5444 5343
rect 6228 5337 6259 5343
rect 7085 5337 7107 5343
rect 7149 5337 7164 5343
rect 93 5317 108 5323
rect 189 5317 204 5323
rect 324 5317 339 5323
rect 445 5317 460 5323
rect 685 5317 723 5323
rect 269 5297 291 5303
rect 717 5297 723 5317
rect 772 5317 787 5323
rect 1293 5317 1315 5323
rect 1373 5317 1395 5323
rect 1700 5317 1731 5323
rect 1725 5297 1731 5317
rect 1981 5317 2003 5323
rect 2100 5317 2131 5323
rect 3197 5317 3212 5323
rect 3437 5317 3452 5323
rect 3508 5317 3523 5323
rect 4093 5317 4108 5323
rect 4269 5317 4307 5323
rect 1741 5297 1779 5303
rect 4269 5297 4275 5317
rect 4413 5317 4492 5323
rect 4804 5317 4819 5323
rect 5037 5317 5075 5323
rect 5037 5297 5043 5317
rect 5204 5317 5219 5323
rect 5501 5317 5516 5323
rect 5645 5317 5683 5323
rect 5316 5296 5324 5304
rect 5677 5297 5683 5317
rect 6509 5317 6547 5323
rect 6541 5297 6547 5317
rect 7085 5324 7091 5337
rect 7108 5317 7123 5323
rect 7149 5317 7187 5323
rect 7149 5297 7155 5317
rect 7316 5317 7331 5323
rect 1389 5277 1484 5283
rect 5092 5277 5107 5283
rect 6570 5276 6572 5284
rect 746 5256 748 5264
rect 1690 5256 1692 5264
rect 858 5236 860 5244
rect 4378 5236 4380 5244
rect 4538 5236 4540 5244
rect 1434 5214 1446 5216
rect 4442 5214 4454 5216
rect 1419 5206 1421 5214
rect 1429 5206 1431 5214
rect 1439 5206 1441 5214
rect 1449 5206 1451 5214
rect 1459 5206 1461 5214
rect 4427 5206 4429 5214
rect 4437 5206 4439 5214
rect 4447 5206 4449 5214
rect 4457 5206 4459 5214
rect 4467 5206 4469 5214
rect 1434 5204 1446 5206
rect 4442 5204 4454 5206
rect 5028 5176 5030 5184
rect 3892 5136 3898 5144
rect 5306 5136 5308 5144
rect 5892 5136 5894 5144
rect 6340 5136 6346 5144
rect 6644 5136 6650 5144
rect 6836 5136 6842 5144
rect 253 5117 275 5123
rect 308 5117 323 5123
rect 644 5117 659 5123
rect 1997 5117 2019 5123
rect 2797 5117 2835 5123
rect 285 5097 300 5103
rect 948 5097 963 5103
rect 1156 5097 1187 5103
rect 1197 5097 1212 5103
rect 1268 5097 1283 5103
rect 1709 5097 1747 5103
rect 2116 5097 2131 5103
rect 2164 5097 2195 5103
rect 2349 5097 2403 5103
rect 2588 5103 2596 5106
rect 2484 5097 2499 5103
rect 2573 5097 2596 5103
rect 2836 5097 2851 5103
rect 3156 5097 3171 5103
rect 3492 5097 3507 5103
rect 4285 5103 4291 5123
rect 4644 5116 4652 5124
rect 4285 5097 4323 5103
rect 4653 5097 4684 5103
rect 4829 5097 4860 5103
rect 4941 5097 4956 5103
rect 4973 5097 5027 5103
rect 5085 5103 5091 5123
rect 5068 5097 5091 5103
rect 5068 5092 5076 5097
rect 5252 5097 5283 5103
rect 5549 5103 5555 5123
rect 5917 5117 5932 5123
rect 7341 5117 7356 5123
rect 5508 5097 5523 5103
rect 5549 5097 5572 5103
rect 5564 5092 5572 5097
rect 5613 5097 5667 5103
rect 5677 5097 5692 5103
rect 5796 5097 5811 5103
rect 6061 5097 6108 5103
rect 573 5077 604 5083
rect 836 5077 851 5083
rect 1133 5077 1148 5083
rect 1533 5077 1571 5083
rect 1677 5077 1692 5083
rect 4028 5077 4052 5083
rect 4900 5077 4931 5083
rect 5245 5077 5267 5083
rect 5492 5077 5507 5083
rect 6205 5077 6243 5083
rect 424 5056 428 5064
rect 1581 5057 1596 5063
rect 3485 5057 3507 5063
rect 5732 5057 5747 5063
rect 6036 5056 6038 5064
rect 6237 5057 6243 5077
rect 6509 5057 6547 5063
rect 7197 5057 7235 5063
rect 360 5036 364 5044
rect 1946 5036 1948 5044
rect 2026 5036 2028 5044
rect 2938 5014 2950 5016
rect 5946 5014 5958 5016
rect 2923 5006 2925 5014
rect 2933 5006 2935 5014
rect 2943 5006 2945 5014
rect 2953 5006 2955 5014
rect 2963 5006 2965 5014
rect 5931 5006 5933 5014
rect 5941 5006 5943 5014
rect 5951 5006 5953 5014
rect 5961 5006 5963 5014
rect 5971 5006 5973 5014
rect 2938 5004 2950 5006
rect 5946 5004 5958 5006
rect 72 4976 76 4984
rect 1492 4977 1507 4983
rect 2644 4976 2646 4984
rect 2996 4977 3011 4983
rect 445 4957 472 4963
rect 692 4957 707 4963
rect 3229 4957 3251 4963
rect 3357 4957 3379 4963
rect 3629 4957 3651 4963
rect 4381 4957 4419 4963
rect 109 4924 115 4943
rect 260 4937 275 4943
rect 820 4937 835 4943
rect 1204 4937 1219 4943
rect 1236 4937 1251 4943
rect 1421 4937 1507 4943
rect 1773 4937 1795 4943
rect 2004 4937 2024 4943
rect 2173 4937 2188 4943
rect 2349 4937 2403 4943
rect 3060 4937 3075 4943
rect 3300 4937 3315 4943
rect 4452 4937 4515 4943
rect 5085 4943 5091 4963
rect 6573 4957 6588 4963
rect 6893 4957 6908 4963
rect 5053 4937 5091 4943
rect 5709 4937 5724 4943
rect 6468 4937 6483 4943
rect 6589 4937 6620 4943
rect 116 4917 140 4923
rect 525 4917 563 4923
rect 925 4917 940 4923
rect 1405 4917 1436 4923
rect 1549 4917 1571 4923
rect 1629 4917 1651 4923
rect 1693 4917 1731 4923
rect 1933 4917 1971 4923
rect 2180 4917 2195 4923
rect 2397 4917 2412 4923
rect 2445 4917 2460 4923
rect 2524 4923 2532 4928
rect 2524 4917 2547 4923
rect 2052 4897 2067 4903
rect 2148 4896 2156 4904
rect 2484 4896 2492 4904
rect 2541 4897 2547 4917
rect 2909 4917 3011 4923
rect 2653 4897 2675 4903
rect 3005 4897 3011 4917
rect 3293 4917 3308 4923
rect 3588 4917 3603 4923
rect 4525 4917 4563 4923
rect 4589 4917 4604 4923
rect 3117 4897 3155 4903
rect 4557 4897 4563 4917
rect 4628 4917 4643 4923
rect 4692 4917 4707 4923
rect 4756 4917 4771 4923
rect 5076 4917 5091 4923
rect 5565 4917 5580 4923
rect 5725 4917 5740 4923
rect 5972 4917 5987 4923
rect 5997 4917 6051 4923
rect 6125 4917 6179 4923
rect 6220 4923 6228 4928
rect 6220 4917 6243 4923
rect 5778 4896 5788 4904
rect 6237 4897 6243 4917
rect 6308 4917 6323 4923
rect 6589 4917 6595 4937
rect 6957 4943 6963 4963
rect 6893 4937 6915 4943
rect 6925 4937 6963 4943
rect 6909 4917 6915 4937
rect 7069 4943 7075 4963
rect 6996 4937 7027 4943
rect 7037 4937 7075 4943
rect 7021 4917 7027 4937
rect 2436 4876 2438 4884
rect 2877 4877 2892 4883
rect 6266 4876 6268 4884
rect 234 4836 236 4844
rect 426 4836 428 4844
rect 794 4836 796 4844
rect 1866 4836 1868 4844
rect 1978 4836 1980 4844
rect 2202 4836 2204 4844
rect 6052 4836 6054 4844
rect 6708 4836 6710 4844
rect 6804 4836 6806 4844
rect 1434 4814 1446 4816
rect 4442 4814 4454 4816
rect 1419 4806 1421 4814
rect 1429 4806 1431 4814
rect 1439 4806 1441 4814
rect 1449 4806 1451 4814
rect 1459 4806 1461 4814
rect 4427 4806 4429 4814
rect 4437 4806 4439 4814
rect 4447 4806 4449 4814
rect 4457 4806 4459 4814
rect 4467 4806 4469 4814
rect 1434 4804 1446 4806
rect 4442 4804 4454 4806
rect 5140 4756 5142 4764
rect 6116 4756 6118 4764
rect 1124 4736 1126 4744
rect 2202 4736 2204 4744
rect 5220 4736 5222 4744
rect 749 4717 771 4723
rect 829 4717 851 4723
rect 1149 4717 1171 4723
rect 1293 4704 1299 4723
rect 77 4697 115 4703
rect 237 4697 252 4703
rect 269 4697 284 4703
rect 61 4677 83 4683
rect 317 4683 323 4703
rect 388 4697 403 4703
rect 685 4697 707 4703
rect 852 4697 867 4703
rect 900 4697 915 4703
rect 1012 4697 1027 4703
rect 1108 4697 1123 4703
rect 1165 4697 1203 4703
rect 1300 4697 1331 4703
rect 1688 4697 1724 4703
rect 1821 4703 1827 4723
rect 3021 4717 3043 4723
rect 3101 4717 3123 4723
rect 4244 4717 4259 4723
rect 4660 4716 4668 4724
rect 1821 4697 1875 4703
rect 2228 4697 2243 4703
rect 2548 4697 2563 4703
rect 2797 4697 2819 4703
rect 3668 4697 3699 4703
rect 3812 4697 3827 4703
rect 4685 4703 4691 4723
rect 4964 4716 4972 4724
rect 4644 4697 4659 4703
rect 4685 4697 4723 4703
rect 4989 4703 4995 4723
rect 4989 4697 5027 4703
rect 5165 4697 5180 4703
rect 5581 4697 5628 4703
rect 5677 4703 5683 4723
rect 5645 4697 5683 4703
rect 6100 4697 6115 4703
rect 6340 4697 6355 4703
rect 317 4677 355 4683
rect 372 4677 387 4683
rect 397 4677 419 4683
rect 93 4657 108 4663
rect 221 4657 236 4663
rect 301 4657 332 4663
rect 381 4657 387 4677
rect 1085 4677 1100 4683
rect 605 4657 620 4663
rect 1085 4657 1091 4677
rect 1229 4677 1244 4683
rect 1229 4657 1235 4677
rect 1501 4677 1516 4683
rect 1981 4677 1996 4683
rect 2013 4677 2051 4683
rect 2221 4677 2243 4683
rect 2468 4677 2483 4683
rect 2660 4676 2664 4684
rect 2749 4677 2803 4683
rect 2861 4677 2899 4683
rect 2909 4677 2988 4683
rect 2152 4656 2156 4664
rect 2260 4657 2275 4663
rect 2909 4657 2915 4677
rect 3053 4677 3068 4683
rect 3053 4657 3059 4677
rect 3549 4677 3564 4683
rect 5597 4677 5612 4683
rect 6461 4677 6476 4683
rect 4588 4664 4596 4672
rect 4109 4657 4131 4663
rect 6036 4657 6051 4663
rect 6477 4657 6483 4676
rect 6493 4657 6531 4663
rect 490 4636 492 4644
rect 1482 4636 1484 4644
rect 3092 4636 3094 4644
rect 3332 4636 3336 4644
rect 2938 4614 2950 4616
rect 5946 4614 5958 4616
rect 2923 4606 2925 4614
rect 2933 4606 2935 4614
rect 2943 4606 2945 4614
rect 2953 4606 2955 4614
rect 2963 4606 2965 4614
rect 5931 4606 5933 4614
rect 5941 4606 5943 4614
rect 5951 4606 5953 4614
rect 5961 4606 5963 4614
rect 5971 4606 5973 4614
rect 2938 4604 2950 4606
rect 5946 4604 5958 4606
rect 264 4576 268 4584
rect 1924 4576 1926 4584
rect 2106 4576 2108 4584
rect 2650 4576 2652 4584
rect 5268 4576 5270 4584
rect 772 4557 803 4563
rect 1140 4556 1148 4564
rect 61 4517 92 4523
rect 205 4523 211 4543
rect 525 4537 547 4543
rect 1629 4537 1651 4543
rect 1693 4537 1715 4543
rect 1940 4537 1955 4543
rect 2045 4537 2060 4543
rect 2525 4537 2540 4543
rect 2845 4537 2883 4543
rect 3114 4536 3116 4544
rect 3629 4537 3644 4543
rect 3908 4537 3923 4543
rect 4525 4543 4531 4563
rect 5485 4557 5523 4563
rect 6045 4557 6060 4563
rect 6765 4557 6803 4563
rect 6877 4557 6915 4563
rect 7005 4557 7028 4563
rect 7020 4554 7028 4557
rect 4493 4537 4531 4543
rect 4989 4537 5011 4543
rect 5060 4537 5075 4543
rect 6733 4537 6748 4543
rect 6948 4537 6979 4543
rect 173 4517 211 4523
rect 381 4517 419 4523
rect 381 4497 387 4517
rect 628 4517 659 4523
rect 717 4517 739 4523
rect 772 4517 787 4523
rect 1092 4517 1107 4523
rect 1421 4517 1468 4523
rect 1549 4517 1587 4523
rect 1716 4517 1731 4523
rect 1805 4517 1820 4523
rect 2068 4517 2083 4523
rect 2557 4517 2572 4523
rect 2932 4517 2979 4523
rect 3741 4517 3779 4523
rect 3821 4517 3859 4523
rect 3885 4517 3916 4523
rect 1540 4496 1548 4504
rect 1885 4497 1900 4503
rect 2077 4497 2099 4503
rect 3853 4497 3859 4517
rect 4420 4517 4476 4523
rect 4573 4517 4588 4523
rect 4652 4523 4660 4528
rect 4637 4517 4660 4523
rect 3965 4497 4003 4503
rect 4637 4497 4643 4517
rect 4973 4517 4988 4523
rect 5197 4517 5212 4523
rect 5293 4517 5308 4523
rect 5645 4517 5660 4523
rect 6308 4517 6323 4523
rect 6372 4517 6387 4523
rect 6428 4523 6436 4528
rect 6428 4517 6451 4523
rect 6445 4497 6451 4517
rect 6973 4517 6979 4537
rect 7341 4537 7404 4543
rect 6989 4517 7004 4523
rect 7085 4517 7100 4523
rect 6090 4456 6092 4464
rect 122 4436 124 4444
rect 602 4436 604 4444
rect 746 4436 748 4444
rect 2436 4436 2438 4444
rect 2804 4436 2806 4444
rect 5092 4436 5094 4444
rect 5172 4436 5174 4444
rect 5412 4436 5414 4444
rect 5620 4436 5622 4444
rect 5901 4437 5916 4443
rect 1434 4414 1446 4416
rect 4442 4414 4454 4416
rect 1419 4406 1421 4414
rect 1429 4406 1431 4414
rect 1439 4406 1441 4414
rect 1449 4406 1451 4414
rect 1459 4406 1461 4414
rect 4427 4406 4429 4414
rect 4437 4406 4439 4414
rect 4447 4406 4449 4414
rect 4457 4406 4459 4414
rect 4467 4406 4469 4414
rect 1434 4404 1446 4406
rect 4442 4404 4454 4406
rect 2260 4376 2262 4384
rect 3508 4376 3510 4384
rect 3620 4376 3622 4384
rect 4762 4376 4764 4384
rect 6244 4356 6246 4364
rect 6701 4337 6716 4343
rect 333 4317 371 4323
rect 445 4317 467 4323
rect 285 4297 307 4303
rect 372 4297 387 4303
rect 756 4297 771 4303
rect 61 4277 83 4283
rect 180 4277 195 4283
rect 717 4277 739 4283
rect 765 4277 771 4297
rect 868 4297 892 4303
rect 932 4297 947 4303
rect 1037 4303 1043 4323
rect 1037 4297 1075 4303
rect 1165 4297 1180 4303
rect 1357 4297 1372 4303
rect 1581 4303 1587 4323
rect 1549 4297 1587 4303
rect 1620 4297 1635 4303
rect 1773 4303 1779 4323
rect 3652 4317 3667 4323
rect 1773 4297 1788 4303
rect 1965 4297 1980 4303
rect 2557 4297 2572 4303
rect 4493 4297 4508 4303
rect 4685 4297 4732 4303
rect 4900 4297 4915 4303
rect 4989 4297 5004 4303
rect 5620 4297 5635 4303
rect 1101 4277 1123 4283
rect 1245 4277 1267 4283
rect 1508 4277 1523 4283
rect 1613 4277 1628 4283
rect 2109 4277 2136 4283
rect 2516 4277 2531 4283
rect 3341 4277 3363 4283
rect 4925 4277 4956 4283
rect 4996 4277 5027 4283
rect 5165 4277 5180 4283
rect 148 4256 156 4264
rect 212 4256 220 4264
rect 1885 4257 1907 4263
rect 2344 4256 2348 4264
rect 2756 4257 2771 4263
rect 4948 4257 4963 4263
rect 5629 4257 5635 4297
rect 5661 4283 5667 4303
rect 5853 4303 5859 4323
rect 5821 4297 5859 4303
rect 6189 4297 6243 4303
rect 6301 4303 6307 4323
rect 6284 4297 6307 4303
rect 6284 4292 6292 4297
rect 6605 4303 6611 4323
rect 6573 4297 6611 4303
rect 6765 4303 6771 4323
rect 6733 4297 6771 4303
rect 6877 4303 6883 4323
rect 6804 4297 6851 4303
rect 6877 4297 6915 4303
rect 7165 4297 7180 4303
rect 5661 4277 5683 4283
rect 6596 4277 6611 4283
rect 548 4236 552 4244
rect 824 4236 828 4244
rect 1764 4236 1766 4244
rect 2090 4236 2092 4244
rect 2500 4236 2502 4244
rect 2938 4214 2950 4216
rect 5946 4214 5958 4216
rect 2923 4206 2925 4214
rect 2933 4206 2935 4214
rect 2943 4206 2945 4214
rect 2953 4206 2955 4214
rect 2963 4206 2965 4214
rect 5931 4206 5933 4214
rect 5941 4206 5943 4214
rect 5951 4206 5953 4214
rect 5961 4206 5963 4214
rect 5971 4206 5973 4214
rect 2938 4204 2950 4206
rect 5946 4204 5958 4206
rect 468 4176 472 4184
rect 696 4176 700 4184
rect 1636 4176 1640 4184
rect 2298 4176 2300 4184
rect 2458 4176 2460 4184
rect 2890 4176 2892 4184
rect 3258 4176 3260 4184
rect 93 4143 99 4163
rect 557 4157 579 4163
rect 845 4157 860 4163
rect 1357 4157 1372 4163
rect 1885 4157 1907 4163
rect 2228 4156 2236 4164
rect 3501 4157 3523 4163
rect 4141 4157 4163 4163
rect 4525 4157 4563 4163
rect 93 4137 108 4143
rect 381 4143 387 4156
rect 173 4137 195 4143
rect 301 4137 323 4143
rect 349 4137 387 4143
rect 740 4137 755 4143
rect 941 4143 947 4156
rect 877 4137 915 4143
rect 941 4137 963 4143
rect 1565 4137 1580 4143
rect 1693 4137 1708 4143
rect 1805 4137 1843 4143
rect 2109 4143 2115 4156
rect 4060 4144 4068 4148
rect 2109 4137 2131 4143
rect 2173 4137 2211 4143
rect 2484 4137 2499 4143
rect 2669 4137 2691 4143
rect 941 4117 956 4123
rect 989 4117 1020 4123
rect 1245 4117 1299 4123
rect 1485 4117 1523 4123
rect 1700 4117 1763 4123
rect 1789 4117 1804 4123
rect 1757 4097 1763 4117
rect 1860 4117 1875 4123
rect 2093 4117 2124 4123
rect 2317 4123 2323 4136
rect 2669 4124 2675 4137
rect 2836 4137 2867 4143
rect 2317 4117 2339 4123
rect 2717 4117 2748 4123
rect 2157 4097 2179 4103
rect 2717 4097 2723 4117
rect 3197 4123 3203 4143
rect 3277 4137 3292 4143
rect 3396 4137 3411 4143
rect 3524 4137 3539 4143
rect 3556 4137 3587 4143
rect 3661 4137 3676 4143
rect 3732 4137 3763 4143
rect 3773 4137 3795 4143
rect 4941 4143 4947 4163
rect 6820 4156 6822 4164
rect 4909 4137 4947 4143
rect 5757 4137 5772 4143
rect 5949 4137 6012 4143
rect 3149 4117 3203 4123
rect 3309 4117 3347 4123
rect 2861 4097 2883 4103
rect 3341 4097 3347 4117
rect 3965 4117 3996 4123
rect 4381 4117 4476 4123
rect 4797 4117 4835 4123
rect 4829 4097 4835 4117
rect 5645 4117 5683 4123
rect 5645 4097 5651 4117
rect 5780 4117 5795 4123
rect 5884 4123 5892 4128
rect 5884 4117 5907 4123
rect 5901 4097 5907 4117
rect 6140 4123 6148 4128
rect 6140 4117 6163 4123
rect 6157 4097 6163 4117
rect 6285 4117 6339 4123
rect 6493 4117 6531 4123
rect 6525 4097 6531 4117
rect 6845 4117 6892 4123
rect 7037 4117 7052 4123
rect 7268 4117 7283 4123
rect 6548 4096 6556 4104
rect 541 4077 556 4083
rect 1124 4077 1139 4083
rect 2580 4077 2595 4083
rect 5620 4056 5622 4064
rect 6100 4056 6102 4064
rect 282 4036 284 4044
rect 404 4036 406 4044
rect 1434 4014 1446 4016
rect 4442 4014 4454 4016
rect 1419 4006 1421 4014
rect 1429 4006 1431 4014
rect 1439 4006 1441 4014
rect 1449 4006 1451 4014
rect 1459 4006 1461 4014
rect 4427 4006 4429 4014
rect 4437 4006 4439 4014
rect 4447 4006 4449 4014
rect 4457 4006 4459 4014
rect 4467 4006 4469 4014
rect 1434 4004 1446 4006
rect 4442 4004 4454 4006
rect 90 3976 92 3984
rect 3956 3976 3958 3984
rect 6692 3956 6694 3964
rect 4324 3936 4330 3944
rect 5124 3936 5126 3944
rect 5258 3936 5260 3944
rect 6388 3936 6390 3944
rect 7133 3937 7148 3943
rect 7236 3936 7242 3944
rect 580 3917 595 3923
rect 820 3917 835 3923
rect 541 3903 547 3916
rect 781 3903 787 3916
rect 468 3897 499 3903
rect 509 3897 547 3903
rect 765 3897 787 3903
rect 1165 3897 1180 3903
rect 1773 3897 1795 3903
rect 2093 3897 2115 3903
rect 2429 3903 2435 3923
rect 2724 3917 2739 3923
rect 3421 3917 3443 3923
rect 2429 3897 2467 3903
rect 3316 3897 3395 3903
rect 3901 3897 3955 3903
rect 5021 3897 5036 3903
rect 5149 3897 5203 3903
rect 5773 3903 5779 3923
rect 5876 3916 5884 3924
rect 5741 3897 5779 3903
rect 5885 3897 5923 3903
rect 221 3877 259 3883
rect 724 3877 755 3883
rect 772 3877 803 3883
rect 1268 3877 1299 3883
rect 1412 3877 1475 3883
rect 1709 3877 1747 3883
rect 548 3856 556 3864
rect 660 3856 668 3864
rect 1149 3857 1187 3863
rect 1220 3857 1235 3863
rect 1741 3857 1747 3877
rect 1844 3877 1859 3883
rect 2029 3877 2051 3883
rect 2212 3877 2227 3883
rect 2909 3877 2924 3883
rect 2932 3877 2995 3883
rect 2989 3864 2995 3877
rect 3357 3877 3379 3883
rect 2292 3857 2307 3863
rect 2797 3857 2819 3863
rect 3229 3857 3260 3863
rect 3357 3863 3363 3877
rect 3741 3877 3795 3883
rect 4109 3877 4131 3883
rect 4221 3877 4236 3883
rect 4788 3877 4803 3883
rect 5917 3883 5923 3897
rect 6477 3897 6492 3903
rect 6797 3903 6803 3923
rect 6820 3916 6828 3924
rect 6717 3897 6739 3903
rect 6765 3897 6803 3903
rect 5917 3877 6003 3883
rect 6429 3877 6451 3883
rect 6733 3883 6739 3897
rect 7284 3897 7315 3903
rect 6733 3877 6748 3883
rect 7036 3877 7052 3883
rect 3341 3857 3363 3863
rect 3468 3863 3476 3866
rect 4316 3864 4324 3872
rect 3460 3857 3476 3863
rect 184 3836 188 3844
rect 984 3836 988 3844
rect 1332 3836 1336 3844
rect 1528 3836 1532 3844
rect 1620 3836 1624 3844
rect 2568 3836 2572 3844
rect 3834 3836 3836 3844
rect 4202 3836 4204 3844
rect 5508 3836 5510 3844
rect 6100 3836 6102 3844
rect 2938 3814 2950 3816
rect 5946 3814 5958 3816
rect 2923 3806 2925 3814
rect 2933 3806 2935 3814
rect 2943 3806 2945 3814
rect 2953 3806 2955 3814
rect 2963 3806 2965 3814
rect 5931 3806 5933 3814
rect 5941 3806 5943 3814
rect 5951 3806 5953 3814
rect 5961 3806 5963 3814
rect 5971 3806 5973 3814
rect 2938 3804 2950 3806
rect 5946 3804 5958 3806
rect 3508 3776 3510 3784
rect 4004 3776 4006 3784
rect 4260 3776 4262 3784
rect 5956 3777 6019 3783
rect 77 3743 83 3763
rect 45 3737 83 3743
rect 404 3737 419 3743
rect 525 3737 547 3743
rect 637 3737 659 3743
rect 925 3737 947 3743
rect 1965 3743 1971 3763
rect 2004 3757 2019 3763
rect 2061 3757 2083 3763
rect 2925 3757 3004 3763
rect 3021 3757 3059 3763
rect 3812 3757 3827 3763
rect 4157 3744 4163 3763
rect 1741 3737 1763 3743
rect 1933 3737 1971 3743
rect 2020 3737 2035 3743
rect 2157 3737 2195 3743
rect 2381 3737 2403 3743
rect 2420 3737 2435 3743
rect 3341 3737 3356 3743
rect 4164 3737 4195 3743
rect 4285 3737 4300 3743
rect 4660 3737 4675 3743
rect 5220 3737 5235 3743
rect 5661 3737 5676 3743
rect 6765 3737 6787 3743
rect 140 3723 148 3728
rect 125 3717 148 3723
rect 493 3717 508 3723
rect 701 3717 716 3723
rect 1085 3723 1091 3736
rect 1021 3717 1091 3723
rect 3348 3717 3363 3723
rect 3468 3717 3491 3723
rect 3468 3712 3476 3717
rect 3789 3717 3804 3723
rect 4957 3717 4995 3723
rect 436 3697 451 3703
rect 3604 3697 3619 3703
rect 4484 3697 4531 3703
rect 4957 3697 4963 3717
rect 5085 3717 5139 3723
rect 5197 3717 5228 3723
rect 5348 3717 5363 3723
rect 5629 3717 5644 3723
rect 5677 3717 5708 3723
rect 5677 3697 5683 3717
rect 6045 3717 6060 3723
rect 6525 3717 6579 3723
rect 6685 3717 6716 3723
rect 7060 3717 7075 3723
rect 6628 3696 6636 3704
rect 1213 3677 1276 3683
rect 1284 3677 1299 3683
rect 1332 3677 1347 3683
rect 2084 3677 2099 3683
rect 2520 3676 2524 3684
rect 3076 3676 3078 3684
rect 3597 3677 3612 3683
rect 3597 3657 3603 3677
rect 5364 3676 5366 3684
rect 6154 3676 6156 3684
rect 6804 3656 6806 3664
rect 7076 3656 7078 3664
rect 344 3636 348 3644
rect 586 3636 588 3644
rect 676 3636 678 3644
rect 1405 3637 1468 3643
rect 2680 3636 2684 3644
rect 6996 3636 6998 3644
rect 7140 3636 7142 3644
rect 1434 3614 1446 3616
rect 4442 3614 4454 3616
rect 1419 3606 1421 3614
rect 1429 3606 1431 3614
rect 1439 3606 1441 3614
rect 1449 3606 1451 3614
rect 1459 3606 1461 3614
rect 4427 3606 4429 3614
rect 4437 3606 4439 3614
rect 4447 3606 4449 3614
rect 4457 3606 4459 3614
rect 4467 3606 4469 3614
rect 1434 3604 1446 3606
rect 4442 3604 4454 3606
rect 1050 3576 1052 3584
rect 4986 3576 4988 3584
rect 5370 3576 5372 3584
rect 6010 3576 6012 3584
rect 3828 3556 3830 3564
rect 2372 3536 2374 3544
rect 4100 3537 4115 3543
rect 733 3517 748 3523
rect 205 3497 220 3503
rect 29 3477 51 3483
rect 141 3477 163 3483
rect 253 3477 275 3483
rect 333 3477 355 3483
rect 436 3477 451 3483
rect 733 3477 739 3517
rect 1348 3517 1363 3523
rect 1837 3517 1875 3523
rect 2084 3516 2092 3524
rect 3341 3517 3363 3523
rect 957 3497 972 3503
rect 1421 3497 1484 3503
rect 1636 3497 1651 3503
rect 2740 3497 2755 3503
rect 1837 3477 1859 3483
rect 1965 3477 1987 3483
rect 2125 3477 2147 3483
rect 2205 3477 2220 3483
rect 2413 3477 2435 3483
rect 2628 3477 2643 3483
rect 2749 3477 2755 3497
rect 3229 3497 3308 3503
rect 3453 3497 3468 3503
rect 3549 3497 3564 3503
rect 3748 3497 3763 3503
rect 3773 3497 3827 3503
rect 4109 3497 4115 3537
rect 4180 3536 4182 3544
rect 4810 3536 4812 3544
rect 4781 3503 4787 3523
rect 4749 3497 4787 3503
rect 4909 3497 4924 3503
rect 4932 3497 4963 3503
rect 5044 3497 5059 3503
rect 5197 3497 5212 3503
rect 5869 3497 5900 3503
rect 5908 3497 5987 3503
rect 6653 3503 6659 3523
rect 6621 3497 6659 3503
rect 6797 3497 6812 3503
rect 7028 3497 7043 3503
rect 2957 3477 3020 3483
rect 3085 3477 3107 3483
rect 3261 3477 3292 3483
rect 1325 3457 1340 3463
rect 2253 3457 2275 3463
rect 714 3436 716 3444
rect 1220 3437 1235 3443
rect 1581 3437 1596 3443
rect 1700 3436 1702 3444
rect 1805 3437 1820 3443
rect 2253 3437 2259 3457
rect 2525 3457 2547 3463
rect 3261 3457 3267 3477
rect 3965 3477 3996 3483
rect 4029 3477 4044 3483
rect 5469 3477 5507 3483
rect 5549 3477 5587 3483
rect 3516 3463 3524 3472
rect 4284 3464 4292 3468
rect 3516 3457 3548 3463
rect 3940 3456 3948 3464
rect 5469 3457 5475 3477
rect 5581 3457 5587 3477
rect 6077 3477 6115 3483
rect 5741 3457 5779 3463
rect 6109 3457 6115 3477
rect 6829 3477 6867 3483
rect 6861 3457 6867 3477
rect 2314 3436 2316 3444
rect 2696 3436 2700 3444
rect 2808 3436 2812 3444
rect 2900 3436 2904 3444
rect 4010 3436 4012 3444
rect 4234 3436 4236 3444
rect 2938 3414 2950 3416
rect 5946 3414 5958 3416
rect 2923 3406 2925 3414
rect 2933 3406 2935 3414
rect 2943 3406 2945 3414
rect 2953 3406 2955 3414
rect 2963 3406 2965 3414
rect 5931 3406 5933 3414
rect 5941 3406 5943 3414
rect 5951 3406 5953 3414
rect 5961 3406 5963 3414
rect 5971 3406 5973 3414
rect 2938 3404 2950 3406
rect 5946 3404 5958 3406
rect 221 3357 243 3363
rect 285 3357 300 3363
rect 317 3357 355 3363
rect 557 3363 563 3383
rect 1389 3377 1452 3383
rect 1613 3377 1628 3383
rect 2701 3377 2723 3383
rect 557 3357 579 3363
rect 2093 3357 2115 3363
rect 2701 3363 2707 3377
rect 2980 3376 2984 3384
rect 3940 3376 3942 3384
rect 2685 3357 2707 3363
rect 3293 3357 3331 3363
rect 4180 3357 4195 3363
rect 5101 3357 5139 3363
rect 6397 3357 6435 3363
rect 29 3337 44 3343
rect 189 3337 211 3343
rect 589 3337 611 3343
rect 2125 3337 2147 3343
rect 2205 3337 2227 3343
rect 2244 3337 2275 3343
rect 2292 3337 2307 3343
rect 2397 3337 2419 3343
rect 2653 3337 2675 3343
rect 2708 3337 2739 3343
rect 4116 3337 4131 3343
rect 4420 3337 4499 3343
rect 7085 3337 7100 3343
rect 61 3317 76 3323
rect 653 3317 668 3323
rect 829 3317 844 3323
rect 1668 3317 1683 3323
rect 1741 3317 1763 3323
rect 1917 3317 1932 3323
rect 2349 3317 2387 3323
rect 148 3296 158 3304
rect 397 3283 403 3303
rect 2349 3297 2355 3317
rect 2740 3317 2755 3323
rect 2820 3317 2835 3323
rect 3620 3317 3635 3323
rect 3900 3317 3923 3323
rect 3900 3314 3908 3317
rect 5021 3317 5059 3323
rect 4292 3297 4307 3303
rect 5021 3297 5027 3317
rect 5629 3317 5667 3323
rect 5629 3297 5635 3317
rect 6100 3317 6115 3323
rect 7044 3317 7059 3323
rect 7085 3317 7123 3323
rect 7085 3297 7091 3317
rect 7316 3317 7331 3323
rect 381 3277 403 3283
rect 445 3277 476 3283
rect 868 3277 899 3283
rect 2020 3277 2051 3283
rect 5878 3276 5884 3284
rect 548 3236 550 3244
rect 1434 3214 1446 3216
rect 4442 3214 4454 3216
rect 1419 3206 1421 3214
rect 1429 3206 1431 3214
rect 1439 3206 1441 3214
rect 1449 3206 1451 3214
rect 1459 3206 1461 3214
rect 4427 3206 4429 3214
rect 4437 3206 4439 3214
rect 4447 3206 4449 3214
rect 4457 3206 4459 3214
rect 4467 3206 4469 3214
rect 1434 3204 1446 3206
rect 4442 3204 4454 3206
rect 2906 3176 2908 3184
rect 6954 3176 6956 3184
rect 2826 3156 2828 3164
rect 804 3137 835 3143
rect 884 3137 899 3143
rect 1156 3137 1171 3143
rect 1309 3137 1363 3143
rect 1508 3137 1539 3143
rect 1805 3137 1820 3143
rect 1917 3137 1948 3143
rect 2490 3136 2492 3144
rect 2749 3137 2764 3143
rect 3860 3137 3875 3143
rect 5322 3136 5324 3144
rect 93 3103 99 3123
rect 2189 3117 2211 3123
rect 4109 3117 4131 3123
rect 4148 3116 4156 3124
rect 5748 3116 5756 3124
rect 93 3097 131 3103
rect 237 3097 252 3103
rect 493 3097 508 3103
rect 29 3077 51 3083
rect 173 3077 195 3083
rect 333 3077 355 3083
rect 413 3077 435 3083
rect 525 3077 547 3083
rect 605 3077 643 3083
rect 797 3077 803 3108
rect 861 3077 867 3108
rect 1101 3097 1116 3103
rect 973 3077 1004 3083
rect 1053 3077 1068 3083
rect 1076 3077 1091 3083
rect 1501 3077 1507 3108
rect 1565 3077 1571 3108
rect 1629 3077 1635 3108
rect 1693 3077 1699 3108
rect 1757 3077 1763 3108
rect 1821 3077 1827 3108
rect 1933 3077 1939 3108
rect 2077 3083 2083 3108
rect 2045 3077 2083 3083
rect 2253 3077 2259 3108
rect 2317 3083 2323 3108
rect 2317 3077 2355 3083
rect 2397 3083 2403 3103
rect 2461 3097 2483 3103
rect 2621 3097 2659 3103
rect 2884 3097 2899 3103
rect 3469 3097 3491 3103
rect 3556 3097 3571 3103
rect 3684 3097 3699 3103
rect 3933 3097 3948 3103
rect 4413 3097 4476 3103
rect 4596 3097 4611 3103
rect 5133 3103 5139 3116
rect 5076 3097 5091 3103
rect 5101 3097 5139 3103
rect 5245 3097 5292 3103
rect 5421 3097 5436 3103
rect 5549 3097 5603 3103
rect 5757 3097 5772 3103
rect 6084 3097 6099 3103
rect 6260 3097 6275 3103
rect 6333 3103 6339 3123
rect 6548 3116 6556 3124
rect 6316 3097 6339 3103
rect 6316 3092 6324 3097
rect 6493 3097 6547 3103
rect 6605 3103 6611 3123
rect 6893 3117 6931 3123
rect 6588 3097 6611 3103
rect 6588 3092 6596 3097
rect 6788 3097 6803 3103
rect 7156 3097 7171 3103
rect 7348 3097 7363 3103
rect 2397 3077 2419 3083
rect 2596 3077 2611 3083
rect 2685 3077 2707 3083
rect 2845 3077 2867 3083
rect 3069 3077 3107 3083
rect 4333 3077 4364 3083
rect 4749 3077 4764 3083
rect 5437 3077 5452 3083
rect 5620 3077 5635 3083
rect 5773 3077 5796 3083
rect 5788 3072 5796 3077
rect 6132 3077 6163 3083
rect 7300 3077 7331 3083
rect 7348 3077 7379 3083
rect 3900 3064 3908 3072
rect 493 3057 515 3063
rect 493 3037 499 3057
rect 2877 3057 2899 3063
rect 2925 3057 2972 3063
rect 676 3036 678 3044
rect 1156 3037 1171 3043
rect 2749 3037 2764 3043
rect 2893 3037 2899 3057
rect 4765 3057 4803 3063
rect 6685 3057 6723 3063
rect 7293 3057 7308 3063
rect 7341 3057 7356 3063
rect 3156 3036 3160 3044
rect 2938 3014 2950 3016
rect 5946 3014 5958 3016
rect 2923 3006 2925 3014
rect 2933 3006 2935 3014
rect 2943 3006 2945 3014
rect 2953 3006 2955 3014
rect 2963 3006 2965 3014
rect 5931 3006 5933 3014
rect 5941 3006 5943 3014
rect 5951 3006 5953 3014
rect 5961 3006 5963 3014
rect 5971 3006 5973 3014
rect 2938 3004 2950 3006
rect 5946 3004 5958 3006
rect 1268 2977 1283 2983
rect 1332 2976 1334 2984
rect 1860 2976 1862 2984
rect 2026 2976 2028 2984
rect 2106 2976 2108 2984
rect 3700 2976 3702 2984
rect 4394 2976 4396 2984
rect 333 2957 355 2963
rect 612 2957 627 2963
rect 701 2957 723 2963
rect 29 2937 51 2943
rect 221 2937 243 2943
rect 301 2937 323 2943
rect 532 2937 547 2943
rect 733 2937 755 2943
rect 797 2937 812 2943
rect 973 2937 995 2943
rect 1053 2937 1075 2943
rect 1181 2937 1196 2943
rect 93 2917 131 2923
rect 93 2897 99 2917
rect 173 2917 204 2923
rect 644 2917 659 2923
rect 797 2917 835 2923
rect 797 2897 803 2917
rect 1037 2917 1052 2923
rect 1092 2917 1123 2923
rect 1245 2912 1251 2943
rect 1581 2937 1635 2943
rect 1821 2937 1843 2943
rect 1885 2943 1891 2963
rect 3412 2957 3427 2963
rect 4276 2957 4291 2963
rect 1876 2937 1891 2943
rect 1965 2937 2003 2943
rect 2052 2937 2083 2943
rect 2253 2937 2291 2943
rect 2349 2937 2371 2943
rect 2509 2937 2531 2943
rect 2589 2937 2611 2943
rect 2948 2937 3011 2943
rect 3373 2937 3443 2943
rect 3725 2937 3756 2943
rect 4060 2943 4068 2944
rect 4060 2937 4076 2943
rect 4324 2937 4355 2943
rect 4637 2937 4675 2943
rect 5277 2943 5283 2963
rect 5277 2937 5315 2943
rect 5389 2937 5404 2943
rect 5869 2943 5875 2956
rect 5869 2937 5891 2943
rect 5988 2937 6019 2943
rect 2148 2917 2163 2923
rect 2173 2917 2211 2923
rect 2573 2917 2588 2923
rect 3972 2917 4003 2923
rect 4253 2917 4284 2923
rect 4436 2917 4499 2923
rect 5348 2917 5363 2923
rect 5389 2917 5427 2923
rect 2676 2897 2691 2903
rect 4644 2897 4659 2903
rect 5389 2897 5395 2917
rect 5892 2917 5907 2923
rect 6676 2917 6691 2923
rect 6749 2917 6788 2923
rect 6780 2914 6788 2917
rect 7124 2917 7139 2923
rect 7284 2917 7299 2923
rect 5908 2896 5916 2904
rect 436 2876 438 2884
rect 1117 2877 1132 2883
rect 2797 2877 2812 2883
rect 2925 2837 2940 2843
rect 6036 2836 6038 2844
rect 6538 2836 6540 2844
rect 6724 2836 6726 2844
rect 1434 2814 1446 2816
rect 4442 2814 4454 2816
rect 1419 2806 1421 2814
rect 1429 2806 1431 2814
rect 1439 2806 1441 2814
rect 1449 2806 1451 2814
rect 1459 2806 1461 2814
rect 4427 2806 4429 2814
rect 4437 2806 4439 2814
rect 4447 2806 4449 2814
rect 4457 2806 4459 2814
rect 4467 2806 4469 2814
rect 1434 2804 1446 2806
rect 4442 2804 4454 2806
rect 2788 2776 2790 2784
rect 6090 2776 6092 2784
rect 509 2743 515 2763
rect 477 2737 515 2743
rect 93 2703 99 2723
rect 477 2717 483 2737
rect 980 2737 995 2743
rect 2858 2736 2860 2744
rect 3908 2737 3939 2743
rect 4556 2732 4564 2736
rect 957 2717 972 2723
rect 1005 2717 1020 2723
rect 1053 2717 1068 2723
rect 1933 2717 1964 2723
rect 4221 2717 4259 2723
rect 5156 2716 5164 2724
rect 6212 2716 6222 2724
rect 93 2697 131 2703
rect 29 2677 51 2683
rect 173 2677 195 2683
rect 253 2677 275 2683
rect 356 2677 371 2683
rect 493 2677 499 2708
rect 637 2677 659 2683
rect 717 2677 739 2683
rect 765 2677 771 2708
rect 1012 2697 1043 2703
rect 1245 2703 1251 2716
rect 1204 2697 1219 2703
rect 1229 2697 1251 2703
rect 1661 2697 1676 2703
rect 1693 2697 1708 2703
rect 1844 2697 1891 2703
rect 2317 2697 2332 2703
rect 2868 2697 2915 2703
rect 2925 2697 2988 2703
rect 3085 2697 3100 2703
rect 3629 2697 3683 2703
rect 4237 2697 4252 2703
rect 1012 2677 1027 2683
rect 1101 2677 1123 2683
rect 1389 2677 1436 2683
rect 1981 2677 2003 2683
rect 2061 2677 2083 2683
rect 2253 2677 2275 2683
rect 2333 2677 2355 2683
rect 2884 2677 2899 2683
rect 3220 2677 3235 2683
rect 3268 2677 3299 2683
rect 3364 2677 3384 2683
rect 3944 2677 3987 2683
rect 4020 2677 4051 2683
rect 4237 2677 4243 2697
rect 5949 2697 6060 2703
rect 6237 2697 6252 2703
rect 6349 2697 6364 2703
rect 6573 2703 6579 2723
rect 6596 2716 6604 2724
rect 6541 2697 6579 2703
rect 6941 2703 6947 2723
rect 6964 2716 6972 2724
rect 6909 2697 6947 2703
rect 7092 2697 7123 2703
rect 5517 2677 5548 2683
rect 6468 2677 6483 2683
rect 285 2657 307 2663
rect 301 2637 307 2657
rect 749 2657 771 2663
rect 1412 2657 1475 2663
rect 1821 2657 1836 2663
rect 4397 2657 4460 2663
rect 5533 2657 5571 2663
rect 600 2636 604 2644
rect 1082 2636 1084 2644
rect 1906 2636 1916 2644
rect 3684 2636 3686 2644
rect 4570 2636 4572 2644
rect 4724 2636 4726 2644
rect 6660 2636 6662 2644
rect 2938 2614 2950 2616
rect 5946 2614 5958 2616
rect 2923 2606 2925 2614
rect 2933 2606 2935 2614
rect 2943 2606 2945 2614
rect 2953 2606 2955 2614
rect 2963 2606 2965 2614
rect 5931 2606 5933 2614
rect 5941 2606 5943 2614
rect 5951 2606 5953 2614
rect 5961 2606 5963 2614
rect 5971 2606 5973 2614
rect 2938 2604 2950 2606
rect 5946 2604 5958 2606
rect 1348 2577 1374 2583
rect 1444 2577 1500 2583
rect 1508 2577 1523 2583
rect 1816 2576 1820 2584
rect 2632 2576 2636 2584
rect 2724 2576 2728 2584
rect 3028 2577 3070 2583
rect 3828 2576 3830 2584
rect 4900 2576 4902 2584
rect 4938 2576 4940 2584
rect 5178 2576 5180 2584
rect 477 2557 499 2563
rect 3140 2557 3155 2563
rect 29 2537 51 2543
rect 173 2537 195 2543
rect 285 2537 307 2543
rect 93 2517 131 2523
rect 93 2497 99 2517
rect 237 2517 275 2523
rect 237 2497 243 2517
rect 301 2512 307 2537
rect 365 2512 371 2543
rect 477 2512 483 2543
rect 509 2537 531 2543
rect 573 2537 588 2543
rect 573 2517 611 2523
rect 573 2497 579 2517
rect 781 2512 787 2543
rect 845 2537 867 2543
rect 957 2537 979 2543
rect 1117 2537 1139 2543
rect 845 2512 851 2537
rect 1197 2537 1219 2543
rect 1405 2537 1516 2543
rect 1885 2537 1900 2543
rect 2301 2537 2316 2543
rect 2381 2537 2403 2543
rect 2525 2537 2547 2543
rect 2564 2537 2579 2543
rect 3709 2537 3724 2543
rect 3853 2537 3868 2543
rect 4029 2537 4067 2543
rect 4100 2537 4131 2543
rect 4653 2537 4691 2543
rect 4788 2537 4803 2543
rect 4957 2537 4995 2543
rect 5012 2537 5027 2543
rect 5037 2537 5075 2543
rect 5085 2537 5123 2543
rect 5220 2537 5235 2543
rect 5453 2543 5459 2563
rect 5453 2537 5491 2543
rect 6077 2543 6083 2563
rect 6045 2537 6083 2543
rect 6349 2537 6364 2543
rect 6620 2543 6628 2548
rect 6605 2537 6628 2543
rect 877 2517 915 2523
rect 909 2497 915 2517
rect 941 2517 956 2523
rect 1293 2517 1340 2523
rect 1565 2517 1603 2523
rect 1613 2517 1651 2523
rect 2125 2517 2163 2523
rect 2461 2517 2499 2523
rect 3245 2517 3260 2523
rect 3613 2517 3628 2523
rect 3917 2517 3955 2523
rect 3949 2504 3955 2517
rect 4340 2517 4371 2523
rect 5108 2517 5139 2523
rect 5293 2517 5308 2523
rect 6820 2517 6835 2523
rect 6893 2517 6931 2523
rect 1556 2497 1571 2503
rect 3741 2497 3756 2503
rect 3988 2497 4003 2503
rect 4660 2497 4675 2503
rect 6500 2496 6508 2504
rect 6925 2497 6931 2517
rect 6948 2496 6956 2504
rect 4780 2484 4788 2488
rect 749 2477 780 2483
rect 813 2477 844 2483
rect 996 2477 1011 2483
rect 1252 2477 1267 2483
rect 1914 2476 1916 2484
rect 4589 2477 4604 2483
rect 4589 2457 4595 2477
rect 4972 2483 4980 2488
rect 4964 2477 4980 2483
rect 5052 2484 5060 2488
rect 68 2436 70 2444
rect 650 2436 652 2444
rect 1066 2436 1068 2444
rect 1434 2414 1446 2416
rect 4442 2414 4454 2416
rect 1419 2406 1421 2414
rect 1429 2406 1431 2414
rect 1439 2406 1441 2414
rect 1449 2406 1451 2414
rect 1459 2406 1461 2414
rect 4427 2406 4429 2414
rect 4437 2406 4439 2414
rect 4447 2406 4449 2414
rect 4457 2406 4459 2414
rect 4467 2406 4469 2414
rect 1434 2404 1446 2406
rect 4442 2404 4454 2406
rect 1898 2376 1900 2384
rect 2852 2376 2856 2384
rect 3018 2376 3020 2384
rect 3204 2376 3206 2384
rect 1700 2337 1715 2343
rect 3274 2336 3276 2344
rect 4004 2337 4035 2343
rect 4276 2337 4291 2343
rect 4685 2337 4716 2343
rect 6980 2337 6995 2343
rect 4124 2332 4132 2336
rect 260 2316 268 2324
rect 349 2317 364 2323
rect 1410 2316 1420 2324
rect 2772 2316 2780 2324
rect 2980 2317 2995 2323
rect 3869 2317 3907 2323
rect 4253 2317 4268 2323
rect 5092 2316 5100 2324
rect 5490 2316 5500 2324
rect 6532 2316 6540 2324
rect 244 2297 259 2303
rect 477 2297 492 2303
rect 61 2277 99 2283
rect 157 2277 179 2283
rect 221 2277 243 2283
rect 301 2277 323 2283
rect 461 2277 476 2283
rect 653 2277 668 2283
rect 749 2277 755 2308
rect 772 2277 792 2283
rect 813 2277 819 2308
rect 1668 2297 1683 2303
rect 1188 2277 1203 2283
rect 333 2257 355 2263
rect 1197 2257 1203 2277
rect 1348 2277 1363 2283
rect 1837 2277 1859 2283
rect 1917 2277 1939 2283
rect 2061 2277 2067 2308
rect 2253 2297 2268 2303
rect 2404 2297 2419 2303
rect 2733 2297 2748 2303
rect 3156 2297 3203 2303
rect 3508 2297 3523 2303
rect 4333 2297 4355 2303
rect 5053 2297 5068 2303
rect 5460 2297 5475 2303
rect 6205 2297 6259 2303
rect 6292 2297 6307 2303
rect 6324 2297 6355 2303
rect 2148 2277 2164 2283
rect 2156 2276 2164 2277
rect 2237 2277 2252 2283
rect 2333 2277 2348 2283
rect 2461 2277 2499 2283
rect 3172 2277 3187 2283
rect 4205 2277 4227 2283
rect 4468 2277 4515 2283
rect 5037 2277 5052 2283
rect 5220 2277 5235 2283
rect 5980 2277 6028 2283
rect 6141 2277 6156 2283
rect 6221 2277 6236 2283
rect 6493 2277 6515 2283
rect 1316 2257 1331 2263
rect 1805 2257 1827 2263
rect 836 2237 851 2243
rect 1005 2237 1020 2243
rect 1949 2237 1955 2263
rect 2093 2257 2108 2263
rect 2356 2257 2371 2263
rect 3709 2257 3731 2263
rect 5354 2256 5356 2264
rect 5709 2257 5747 2263
rect 6388 2256 6390 2264
rect 6676 2256 6678 2264
rect 2612 2236 2616 2244
rect 2938 2214 2950 2216
rect 5946 2214 5958 2216
rect 2923 2206 2925 2214
rect 2933 2206 2935 2214
rect 2943 2206 2945 2214
rect 2953 2206 2955 2214
rect 2963 2206 2965 2214
rect 5931 2206 5933 2214
rect 5941 2206 5943 2214
rect 5951 2206 5953 2214
rect 5961 2206 5963 2214
rect 5971 2206 5973 2214
rect 2938 2204 2950 2206
rect 5946 2204 5958 2206
rect 330 2176 332 2184
rect 456 2176 460 2184
rect 554 2176 556 2184
rect 1053 2177 1068 2183
rect 1901 2177 1916 2183
rect 2632 2176 2636 2184
rect 2746 2176 2748 2184
rect 2840 2176 2844 2184
rect 4074 2176 4076 2184
rect 4397 2177 4460 2183
rect 660 2157 675 2163
rect 2701 2157 2716 2163
rect 5133 2157 5171 2163
rect 125 2137 140 2143
rect 168 2136 172 2144
rect 260 2117 291 2123
rect 381 2117 396 2123
rect 605 2117 620 2123
rect 957 2112 963 2143
rect 1021 2112 1027 2143
rect 1085 2112 1091 2143
rect 1149 2112 1155 2143
rect 1364 2137 1379 2143
rect 1252 2117 1267 2123
rect 1565 2112 1571 2143
rect 1741 2112 1747 2143
rect 1805 2112 1811 2143
rect 1933 2137 1971 2143
rect 2013 2137 2035 2143
rect 2013 2117 2019 2137
rect 2260 2137 2275 2143
rect 2285 2123 2291 2143
rect 2349 2137 2364 2143
rect 2477 2123 2483 2143
rect 2285 2117 2307 2123
rect 2429 2117 2483 2123
rect 3101 2123 3107 2143
rect 3588 2137 3603 2143
rect 3821 2137 3836 2143
rect 3869 2137 3891 2143
rect 4164 2137 4179 2143
rect 5012 2137 5027 2143
rect 5629 2143 5635 2163
rect 6701 2157 6739 2163
rect 5597 2137 5635 2143
rect 5988 2137 6019 2143
rect 6420 2137 6435 2143
rect 6468 2137 6483 2143
rect 6724 2137 6755 2143
rect 3021 2117 3075 2123
rect 3101 2117 3160 2123
rect 1124 2077 1171 2083
rect 1549 2083 1555 2103
rect 3069 2097 3075 2117
rect 3316 2117 3347 2123
rect 3357 2117 3395 2123
rect 3453 2117 3507 2123
rect 3757 2117 3788 2123
rect 4509 2117 4531 2123
rect 4845 2117 4876 2123
rect 4989 2117 5027 2123
rect 3293 2097 3331 2103
rect 3853 2097 3868 2103
rect 5021 2097 5027 2117
rect 5076 2117 5091 2123
rect 5309 2117 5324 2123
rect 6253 2117 6268 2123
rect 6413 2117 6428 2123
rect 6445 2117 6483 2123
rect 6477 2097 6483 2117
rect 6829 2117 6867 2123
rect 6861 2097 6867 2117
rect 7229 2117 7244 2123
rect 7268 2117 7283 2123
rect 1549 2077 1587 2083
rect 1444 2057 1507 2063
rect 1581 2057 1587 2077
rect 4918 2076 4924 2084
rect 4957 2077 4972 2083
rect 6326 2076 6332 2084
rect 6413 2077 6428 2083
rect 234 2036 236 2044
rect 1434 2014 1446 2016
rect 4442 2014 4454 2016
rect 1419 2006 1421 2014
rect 1429 2006 1431 2014
rect 1439 2006 1441 2014
rect 1449 2006 1451 2014
rect 1459 2006 1461 2014
rect 4427 2006 4429 2014
rect 4437 2006 4439 2014
rect 4447 2006 4449 2014
rect 4457 2006 4459 2014
rect 4467 2006 4469 2014
rect 1434 2004 1446 2006
rect 4442 2004 4454 2006
rect 564 1976 566 1984
rect 788 1976 790 1984
rect 2196 1976 2198 1984
rect 2244 1976 2246 1984
rect 2676 1976 2680 1984
rect 2772 1976 2774 1984
rect 3364 1976 3366 1984
rect 6132 1976 6134 1984
rect 237 1937 291 1943
rect 909 1937 940 1943
rect 1101 1937 1116 1943
rect 1332 1937 1363 1943
rect 1501 1937 1516 1943
rect 2394 1936 2396 1944
rect 2468 1937 2515 1943
rect 2548 1937 2579 1943
rect 2797 1937 2812 1943
rect 3242 1936 3244 1944
rect 4788 1937 4819 1943
rect 5684 1936 5686 1944
rect 6461 1937 6476 1943
rect 4652 1932 4660 1936
rect 1037 1917 1052 1923
rect 2292 1916 2300 1924
rect 2589 1917 2604 1923
rect 2884 1916 2892 1924
rect 2932 1917 2995 1923
rect 3117 1917 3155 1923
rect 3453 1917 3491 1923
rect 3508 1917 3523 1923
rect 3533 1917 3571 1923
rect 4653 1917 4668 1923
rect 4701 1917 4723 1923
rect 4772 1917 4787 1923
rect 5156 1916 5164 1924
rect 157 1897 172 1903
rect 77 1877 99 1883
rect 157 1877 163 1897
rect 381 1897 396 1903
rect 797 1897 819 1903
rect 1773 1897 1788 1903
rect 2020 1897 2035 1903
rect 2132 1897 2147 1903
rect 2253 1897 2268 1903
rect 2740 1897 2755 1903
rect 733 1877 771 1883
rect 436 1857 451 1863
rect 765 1857 771 1877
rect 1676 1877 1692 1883
rect 1676 1876 1684 1877
rect 1900 1877 1916 1883
rect 1900 1876 1908 1877
rect 2333 1877 2355 1883
rect 1197 1857 1212 1863
rect 1965 1857 1980 1863
rect 2365 1857 2387 1863
rect 237 1837 252 1843
rect 1837 1837 1852 1843
rect 2381 1837 2387 1857
rect 2436 1856 2444 1864
rect 2749 1857 2755 1897
rect 2829 1897 2860 1903
rect 3316 1897 3363 1903
rect 3437 1897 3452 1903
rect 3597 1897 3635 1903
rect 3332 1877 3347 1883
rect 3757 1883 3763 1903
rect 3965 1897 3996 1903
rect 4084 1897 4115 1903
rect 4573 1897 4595 1903
rect 5181 1903 5187 1923
rect 6948 1916 6956 1924
rect 5181 1897 5219 1903
rect 5421 1897 5452 1903
rect 5837 1897 5852 1903
rect 6077 1897 6092 1903
rect 6253 1897 6284 1903
rect 6324 1897 6339 1903
rect 3757 1877 3772 1883
rect 3876 1877 3891 1883
rect 4525 1877 4563 1883
rect 4525 1857 4531 1877
rect 4637 1877 4675 1883
rect 4685 1877 4700 1883
rect 5588 1877 5619 1883
rect 5652 1877 5667 1883
rect 5860 1877 5875 1883
rect 6269 1877 6307 1883
rect 6652 1866 6660 1876
rect 5261 1857 5299 1863
rect 5565 1857 5603 1863
rect 6052 1856 6054 1864
rect 6829 1857 6867 1863
rect 2520 1836 2524 1844
rect 5812 1836 5814 1844
rect 6458 1836 6460 1844
rect 2938 1814 2950 1816
rect 5946 1814 5958 1816
rect 2923 1806 2925 1814
rect 2933 1806 2935 1814
rect 2943 1806 2945 1814
rect 2953 1806 2955 1814
rect 2963 1806 2965 1814
rect 5931 1806 5933 1814
rect 5941 1806 5943 1814
rect 5951 1806 5953 1814
rect 5961 1806 5963 1814
rect 5971 1806 5973 1814
rect 2938 1804 2950 1806
rect 5946 1804 5958 1806
rect 980 1776 984 1784
rect 253 1757 268 1763
rect 548 1757 563 1763
rect 1085 1763 1091 1783
rect 1085 1757 1107 1763
rect 29 1737 51 1743
rect 141 1737 163 1743
rect 221 1737 236 1743
rect 276 1737 291 1743
rect 349 1737 371 1743
rect 493 1737 531 1743
rect 644 1737 659 1743
rect 868 1737 899 1743
rect 1229 1743 1235 1763
rect 1389 1763 1395 1783
rect 1389 1757 1411 1763
rect 1588 1757 1603 1763
rect 1117 1737 1139 1743
rect 1197 1737 1219 1743
rect 1229 1737 1244 1743
rect 1261 1737 1283 1743
rect 1421 1737 1507 1743
rect 1613 1743 1619 1763
rect 1748 1757 1763 1763
rect 1613 1737 1651 1743
rect 1773 1743 1779 1763
rect 2461 1763 2467 1783
rect 2884 1776 2888 1784
rect 3988 1776 3990 1784
rect 4100 1776 4102 1784
rect 2445 1757 2467 1763
rect 1773 1737 1811 1743
rect 2013 1737 2035 1743
rect 2052 1737 2067 1743
rect 2125 1737 2147 1743
rect 2164 1737 2179 1743
rect 2237 1737 2259 1743
rect 2340 1737 2355 1743
rect 2413 1737 2435 1743
rect 2548 1737 2563 1743
rect 2621 1737 2643 1743
rect 2733 1743 2739 1763
rect 2749 1757 2764 1763
rect 3309 1757 3331 1763
rect 3885 1757 3907 1763
rect 4292 1757 4307 1763
rect 2724 1737 2739 1743
rect 4365 1737 4387 1743
rect 269 1717 284 1723
rect 436 1717 451 1723
rect 1725 1717 1747 1723
rect 1933 1717 1948 1723
rect 2068 1717 2083 1723
rect 3053 1717 3076 1723
rect 3068 1714 3076 1717
rect 3581 1717 3596 1723
rect 3812 1717 3859 1723
rect 4157 1717 4179 1723
rect 4269 1717 4291 1723
rect 4301 1717 4339 1723
rect 4413 1717 4476 1723
rect 308 1696 316 1704
rect 1444 1697 1484 1703
rect 2386 1696 2396 1704
rect 2580 1696 2588 1704
rect 4333 1697 4339 1717
rect 4589 1717 4611 1723
rect 4733 1723 4739 1743
rect 4797 1737 4828 1743
rect 4925 1737 4940 1743
rect 6868 1737 6883 1743
rect 7021 1737 7036 1743
rect 4628 1717 4643 1723
rect 4701 1717 4739 1723
rect 4749 1717 4780 1723
rect 4813 1717 4851 1723
rect 4861 1717 4883 1723
rect 5117 1717 5132 1723
rect 4813 1697 4819 1717
rect 5357 1717 5372 1723
rect 5629 1717 5644 1723
rect 6308 1717 6339 1723
rect 6477 1717 6492 1723
rect 6748 1723 6756 1728
rect 6733 1717 6756 1723
rect 5684 1696 5692 1704
rect 6733 1697 6739 1717
rect 6797 1717 6812 1723
rect 7069 1717 7107 1723
rect 7101 1697 7107 1717
rect 7229 1717 7244 1723
rect 7124 1696 7132 1704
rect 1892 1677 1907 1683
rect 3108 1676 3114 1684
rect 3485 1677 3500 1683
rect 5818 1656 5820 1664
rect 2964 1637 3027 1643
rect 4580 1636 4582 1644
rect 5604 1636 5606 1644
rect 6452 1636 6454 1644
rect 6580 1636 6582 1644
rect 1434 1614 1446 1616
rect 4442 1614 4454 1616
rect 1419 1606 1421 1614
rect 1429 1606 1431 1614
rect 1439 1606 1441 1614
rect 1449 1606 1451 1614
rect 1459 1606 1461 1614
rect 4427 1606 4429 1614
rect 4437 1606 4439 1614
rect 4447 1606 4449 1614
rect 4457 1606 4459 1614
rect 4467 1606 4469 1614
rect 1434 1604 1446 1606
rect 4442 1604 4454 1606
rect 1421 1577 1484 1583
rect 1672 1576 1676 1584
rect 2010 1576 2012 1584
rect 2564 1576 2566 1584
rect 6212 1576 6214 1584
rect 692 1537 723 1543
rect 1156 1536 1160 1544
rect 1236 1537 1251 1543
rect 4573 1537 4620 1543
rect 4044 1532 4052 1536
rect 626 1516 636 1524
rect 413 1483 419 1503
rect 493 1497 515 1503
rect 861 1503 867 1523
rect 829 1497 867 1503
rect 989 1497 1011 1503
rect 1021 1497 1036 1503
rect 1572 1497 1587 1503
rect 1981 1497 2003 1503
rect 2084 1497 2099 1503
rect 2413 1497 2428 1503
rect 3044 1497 3059 1503
rect 3181 1497 3196 1503
rect 3549 1503 3555 1523
rect 4237 1517 4259 1523
rect 4596 1517 4611 1523
rect 3508 1497 3523 1503
rect 3549 1497 3587 1503
rect 4173 1497 4211 1503
rect 404 1477 419 1483
rect 477 1477 492 1483
rect 941 1477 972 1483
rect 1725 1483 1731 1496
rect 1709 1477 1731 1483
rect 1885 1477 1900 1483
rect 2676 1477 2691 1483
rect 2765 1477 2787 1483
rect 2765 1464 2771 1477
rect 3428 1477 3459 1483
rect 3764 1477 3779 1483
rect 4205 1477 4211 1497
rect 4973 1497 4988 1503
rect 5197 1497 5212 1503
rect 6237 1497 6252 1503
rect 6541 1497 6556 1503
rect 7005 1503 7011 1523
rect 6973 1497 7011 1503
rect 7117 1497 7132 1503
rect 5149 1477 5187 1483
rect 836 1456 844 1464
rect 932 1457 947 1463
rect 1277 1457 1299 1463
rect 1773 1457 1788 1463
rect 2029 1457 2067 1463
rect 2189 1457 2211 1463
rect 3245 1457 3267 1463
rect 4052 1456 4060 1464
rect 4228 1456 4236 1464
rect 5149 1457 5155 1477
rect 5485 1477 5516 1483
rect 5549 1477 5564 1483
rect 6388 1477 6403 1483
rect 7117 1477 7155 1483
rect 5357 1457 5395 1463
rect 5789 1457 5827 1463
rect 7117 1457 7123 1477
rect 7277 1457 7315 1463
rect 2804 1436 2806 1444
rect 3898 1436 3900 1444
rect 2938 1414 2950 1416
rect 5946 1414 5958 1416
rect 2923 1406 2925 1414
rect 2933 1406 2935 1414
rect 2943 1406 2945 1414
rect 2953 1406 2955 1414
rect 2963 1406 2965 1414
rect 5931 1406 5933 1414
rect 5941 1406 5943 1414
rect 5951 1406 5953 1414
rect 5961 1406 5963 1414
rect 5971 1406 5973 1414
rect 2938 1404 2950 1406
rect 5946 1404 5958 1406
rect 660 1376 662 1384
rect 2520 1376 2524 1384
rect 2941 1377 3004 1383
rect 3956 1377 3971 1383
rect 253 1357 268 1363
rect 1533 1357 1548 1363
rect 1844 1357 1859 1363
rect 1892 1356 1900 1364
rect 2813 1357 2835 1363
rect 3261 1357 3283 1363
rect 45 1337 76 1343
rect 829 1337 844 1343
rect 1197 1337 1212 1343
rect 1341 1343 1347 1356
rect 1245 1337 1283 1343
rect 1341 1337 1363 1343
rect 1540 1337 1571 1343
rect 1757 1337 1779 1343
rect 1917 1337 1955 1343
rect 1965 1337 1996 1343
rect 500 1317 515 1323
rect 669 1317 691 1323
rect 669 1304 675 1317
rect 1165 1317 1180 1323
rect 1389 1317 1491 1323
rect 1965 1317 1971 1337
rect 2157 1343 2163 1356
rect 4252 1352 4260 1356
rect 2036 1337 2067 1343
rect 2141 1337 2163 1343
rect 2237 1337 2275 1343
rect 2084 1317 2099 1323
rect 2461 1323 2467 1343
rect 2612 1337 2643 1343
rect 3332 1337 3347 1343
rect 6157 1337 6179 1343
rect 6228 1337 6243 1343
rect 6285 1337 6307 1343
rect 6420 1337 6451 1343
rect 2461 1317 2492 1323
rect 2669 1317 2691 1323
rect 2772 1317 2787 1323
rect 3725 1317 3763 1323
rect 4125 1317 4147 1323
rect 4845 1317 4883 1323
rect 877 1297 892 1303
rect 1380 1296 1388 1304
rect 4877 1297 4883 1317
rect 5293 1317 5324 1323
rect 5485 1317 5500 1323
rect 6141 1317 6172 1323
rect 6244 1317 6259 1323
rect 6509 1317 6547 1323
rect 4900 1296 4908 1304
rect 6116 1296 6126 1304
rect 6541 1297 6547 1317
rect 6829 1317 6867 1323
rect 6861 1297 6867 1317
rect 6884 1296 6892 1304
rect 3821 1277 3852 1283
rect 3917 1277 3964 1283
rect 6394 1276 6396 1284
rect 1620 1236 1622 1244
rect 3770 1236 3772 1244
rect 5924 1236 5926 1244
rect 6570 1236 6572 1244
rect 1434 1214 1446 1216
rect 4442 1214 4454 1216
rect 1419 1206 1421 1214
rect 1429 1206 1431 1214
rect 1439 1206 1441 1214
rect 1449 1206 1451 1214
rect 1459 1206 1461 1214
rect 4427 1206 4429 1214
rect 4437 1206 4439 1214
rect 4447 1206 4449 1214
rect 4457 1206 4459 1214
rect 4467 1206 4469 1214
rect 1434 1204 1446 1206
rect 4442 1204 4454 1206
rect 202 1176 204 1184
rect 2020 1176 2022 1184
rect 4413 1177 4476 1183
rect 5540 1176 5542 1184
rect 5626 1176 5628 1184
rect 5818 1176 5820 1184
rect 6010 1176 6012 1184
rect 4436 1157 4499 1163
rect 6138 1156 6140 1164
rect 1668 1136 1672 1144
rect 4317 1137 4332 1143
rect 4340 1137 4403 1143
rect 4573 1137 4588 1143
rect 4637 1137 4652 1143
rect 4868 1137 4883 1143
rect 6980 1136 6982 1144
rect 7060 1136 7066 1144
rect 1780 1117 1795 1123
rect 45 1097 67 1103
rect 205 1097 220 1103
rect 61 1084 67 1097
rect 397 1097 419 1103
rect 573 1097 611 1103
rect 621 1097 652 1103
rect 996 1097 1011 1103
rect 1069 1097 1084 1103
rect 1348 1097 1363 1103
rect 1444 1097 1507 1103
rect 2893 1097 2908 1103
rect 3348 1097 3363 1103
rect 3821 1097 3843 1103
rect 5460 1097 5475 1103
rect 5565 1103 5571 1123
rect 5565 1097 5588 1103
rect 5580 1092 5588 1097
rect 5693 1097 5708 1103
rect 5821 1097 5875 1103
rect 6109 1103 6115 1123
rect 6077 1097 6115 1103
rect 6509 1103 6515 1123
rect 6372 1097 6387 1103
rect 6477 1097 6515 1103
rect 6868 1097 6883 1103
rect 7085 1097 7100 1103
rect 7124 1097 7139 1103
rect 461 1077 476 1083
rect 541 1077 579 1083
rect 1133 1077 1187 1083
rect 1213 1077 1251 1083
rect 1341 1077 1356 1083
rect 1213 1057 1219 1077
rect 1524 1077 1555 1083
rect 1828 1077 1852 1083
rect 1885 1077 1907 1083
rect 1901 1064 1907 1077
rect 2468 1077 2483 1083
rect 3485 1077 3500 1083
rect 5140 1077 5156 1083
rect 5732 1077 5747 1083
rect 7196 1077 7212 1083
rect 7268 1077 7283 1083
rect 1380 1056 1388 1064
rect 1860 1056 1868 1064
rect 4164 1057 4188 1063
rect 5117 1057 5132 1063
rect 5389 1057 5427 1063
rect 7229 1057 7267 1063
rect 120 1036 124 1044
rect 458 1036 460 1044
rect 932 1036 934 1044
rect 2932 1037 2995 1043
rect 3898 1036 3900 1044
rect 4042 1036 4044 1044
rect 2938 1014 2950 1016
rect 5946 1014 5958 1016
rect 2923 1006 2925 1014
rect 2933 1006 2935 1014
rect 2943 1006 2945 1014
rect 2953 1006 2955 1014
rect 2963 1006 2965 1014
rect 5931 1006 5933 1014
rect 5941 1006 5943 1014
rect 5951 1006 5953 1014
rect 5961 1006 5963 1014
rect 5971 1006 5973 1014
rect 2938 1004 2950 1006
rect 5946 1004 5958 1006
rect 232 976 236 984
rect 698 976 700 984
rect 794 976 796 984
rect 740 957 755 963
rect 2301 957 2332 963
rect 2413 957 2428 963
rect 3645 957 3667 963
rect 4132 957 4156 963
rect 4637 957 4652 963
rect 948 937 979 943
rect 1613 937 1628 943
rect 2397 937 2451 943
rect 2445 924 2451 937
rect 3114 936 3116 944
rect 3869 937 3900 943
rect 3917 937 3932 943
rect 4029 937 4067 943
rect 4804 937 4819 943
rect 4829 937 4860 943
rect 5556 937 5571 943
rect 5988 937 6003 943
rect 6045 937 6067 943
rect 6317 937 6332 943
rect 7252 937 7267 943
rect 7277 937 7308 943
rect 557 917 572 923
rect 589 917 611 923
rect 676 917 691 923
rect 685 897 691 917
rect 941 917 956 923
rect 989 917 1011 923
rect 1005 904 1011 917
rect 1773 917 1811 923
rect 3709 917 3724 923
rect 4077 917 4092 923
rect 4557 917 4595 923
rect 4701 917 4739 923
rect 4852 917 4867 923
rect 4973 917 5011 923
rect 5028 917 5059 923
rect 5188 917 5203 923
rect 5244 923 5252 928
rect 5244 917 5267 923
rect 5293 917 5308 923
rect 1085 897 1107 903
rect 3741 897 3756 903
rect 3972 897 3987 903
rect 4756 897 4771 903
rect 5261 897 5267 917
rect 5476 917 5491 923
rect 6004 917 6019 923
rect 6196 917 6211 923
rect 6324 917 6355 923
rect 6541 917 6556 923
rect 6684 923 6692 928
rect 6628 917 6643 923
rect 6669 917 6692 923
rect 5492 896 5500 904
rect 6669 897 6675 917
rect 6733 917 6787 923
rect 6877 917 6892 923
rect 6973 917 6988 923
rect 4764 884 4772 888
rect 372 877 387 883
rect 404 877 419 883
rect 1556 876 1560 884
rect 1876 876 1880 884
rect 3268 876 3274 884
rect 4781 877 4796 883
rect 6084 876 6086 884
rect 6708 836 6710 844
rect 6852 836 6854 844
rect 6948 836 6950 844
rect 1434 814 1446 816
rect 4442 814 4454 816
rect 1419 806 1421 814
rect 1429 806 1431 814
rect 1439 806 1441 814
rect 1449 806 1451 814
rect 1459 806 1461 814
rect 4427 806 4429 814
rect 4437 806 4439 814
rect 4447 806 4449 814
rect 4457 806 4459 814
rect 4467 806 4469 814
rect 1434 804 1446 806
rect 4442 804 4454 806
rect 2756 776 2758 784
rect 4020 776 4022 784
rect 4260 776 4262 784
rect 6228 776 6230 784
rect 6612 776 6614 784
rect 6996 776 6998 784
rect 7236 776 7238 784
rect 7364 776 7366 784
rect 324 736 326 744
rect 570 736 572 744
rect 4154 736 4156 744
rect 4820 737 4835 743
rect 1044 717 1059 723
rect 1780 716 1790 724
rect 4084 717 4099 723
rect 5612 706 5620 716
rect 308 697 323 703
rect 509 697 540 703
rect 829 697 844 703
rect 884 697 899 703
rect 1693 697 1715 703
rect 2004 697 2035 703
rect 2196 697 2211 703
rect 2621 697 2659 703
rect 2676 697 2691 703
rect 2829 697 2851 703
rect 4004 697 4019 703
rect 4221 697 4236 703
rect 5101 697 5139 703
rect 5277 697 5315 703
rect 6333 697 6387 703
rect 7197 697 7212 703
rect 7268 697 7283 703
rect 45 677 76 683
rect 140 677 156 683
rect 140 676 148 677
rect 397 677 428 683
rect 372 657 387 663
rect 397 657 403 677
rect 685 677 700 683
rect 724 677 739 683
rect 861 677 915 683
rect 1101 677 1116 683
rect 676 657 691 663
rect 1101 657 1107 677
rect 1325 677 1340 683
rect 1645 677 1683 683
rect 1549 657 1564 663
rect 1645 657 1651 677
rect 2541 677 2579 683
rect 2605 677 2620 683
rect 2653 677 2675 683
rect 2717 677 2739 683
rect 3981 677 4003 683
rect 3228 664 3236 672
rect 3981 664 3987 677
rect 4228 677 4243 683
rect 5876 677 5956 683
rect 6276 677 6291 683
rect 6349 677 6364 683
rect 6404 677 6419 683
rect 6461 677 6476 683
rect 6525 677 6540 683
rect 6653 677 6668 683
rect 7101 677 7139 683
rect 4540 666 4548 676
rect 4924 666 4932 676
rect 2836 657 2851 663
rect 2925 657 2940 663
rect 3437 657 3459 663
rect 3757 657 3779 663
rect 4836 656 4844 664
rect 5821 657 5859 663
rect 5869 657 5932 663
rect 7101 657 7107 677
rect 7156 657 7171 663
rect 7181 657 7196 663
rect 1492 636 1494 644
rect 2938 614 2950 616
rect 5946 614 5958 616
rect 2923 606 2925 614
rect 2933 606 2935 614
rect 2943 606 2945 614
rect 2953 606 2955 614
rect 2963 606 2965 614
rect 5931 606 5933 614
rect 5941 606 5943 614
rect 5951 606 5953 614
rect 5961 606 5963 614
rect 5971 606 5973 614
rect 2938 604 2950 606
rect 5946 604 5958 606
rect 152 576 156 584
rect 1108 576 1112 584
rect 1572 576 1576 584
rect 2468 576 2470 584
rect 20 557 35 563
rect 317 557 355 563
rect 388 556 396 564
rect 452 557 467 563
rect 644 557 668 563
rect 2420 556 2428 564
rect 3101 557 3123 563
rect 5693 557 5731 563
rect 77 543 83 556
rect 77 537 99 543
rect 708 537 739 543
rect 1053 537 1075 543
rect 29 517 44 523
rect 621 523 627 536
rect 1053 524 1059 537
rect 1373 537 1420 543
rect 1716 537 1731 543
rect 1949 543 1955 556
rect 1933 537 1955 543
rect 1988 537 2003 543
rect 2173 537 2188 543
rect 2349 537 2364 543
rect 3612 543 3620 548
rect 3597 537 3620 543
rect 5220 537 5235 543
rect 5357 537 5372 543
rect 5757 537 5788 543
rect 5885 537 5948 543
rect 6388 537 6403 543
rect 605 517 627 523
rect 765 517 819 523
rect 884 517 899 523
rect 1261 523 1267 536
rect 1245 517 1267 523
rect 1412 517 1491 523
rect 1604 517 1651 523
rect 1741 517 1763 523
rect 1853 517 1891 523
rect 1965 517 1987 523
rect 2045 517 2060 523
rect 2077 517 2131 523
rect 2548 517 2579 523
rect 2861 517 2899 523
rect 2925 517 3011 523
rect 3069 517 3091 523
rect 3853 517 3868 523
rect 4324 517 4339 523
rect 4420 517 4483 523
rect 4733 517 4771 523
rect 5133 517 5171 523
rect 5389 517 5427 523
rect 5837 517 5875 523
rect 6365 517 6403 523
rect 420 497 435 503
rect 756 497 771 503
rect 1428 497 1468 503
rect 2381 497 2396 503
rect 6397 497 6403 517
rect 6477 517 6515 523
rect 6509 497 6515 517
rect 6541 517 6556 523
rect 6829 517 6867 523
rect 6861 497 6867 517
rect 6884 496 6892 504
rect 234 476 236 484
rect 2260 477 2275 483
rect 1914 436 1916 444
rect 1434 414 1446 416
rect 4442 414 4454 416
rect 1419 406 1421 414
rect 1429 406 1431 414
rect 1439 406 1441 414
rect 1449 406 1451 414
rect 1459 406 1461 414
rect 4427 406 4429 414
rect 4437 406 4439 414
rect 4447 406 4449 414
rect 4457 406 4459 414
rect 4467 406 4469 414
rect 1434 404 1446 406
rect 4442 404 4454 406
rect 52 376 56 384
rect 148 376 150 384
rect 1754 376 1756 384
rect 7002 376 7004 384
rect 842 336 844 344
rect 954 336 956 344
rect 6740 336 6742 344
rect 173 317 188 323
rect 562 316 572 324
rect 637 317 659 323
rect 1172 316 1180 324
rect 1581 317 1596 323
rect 1645 317 1683 323
rect 1700 317 1731 323
rect 2941 317 3004 323
rect 3076 317 3091 323
rect 3181 317 3203 323
rect 461 297 499 303
rect 852 297 883 303
rect 1028 297 1043 303
rect 1565 297 1580 303
rect 1757 297 1788 303
rect 1796 297 1811 303
rect 1844 297 1859 303
rect 2372 297 2387 303
rect 2397 297 2412 303
rect 2557 297 2579 303
rect 2781 297 2819 303
rect 3156 297 3187 303
rect 3236 297 3251 303
rect 3357 297 3395 303
rect 397 283 403 296
rect 3981 297 4019 303
rect 4685 297 4700 303
rect 5212 303 5220 304
rect 5181 297 5220 303
rect 5581 297 5619 303
rect 5725 297 5740 303
rect 5780 297 5811 303
rect 6204 303 6212 306
rect 6204 297 6227 303
rect 6317 303 6323 323
rect 6317 297 6355 303
rect 6484 297 6499 303
rect 7245 297 7260 303
rect 228 277 259 283
rect 397 277 419 283
rect 516 277 531 283
rect 644 277 659 283
rect 701 277 716 283
rect 1421 277 1532 283
rect 1780 277 1795 283
rect 1837 277 1852 283
rect 1901 277 1955 283
rect 2548 277 2563 283
rect 2621 277 2659 283
rect 2701 277 2739 283
rect 2813 277 2835 283
rect 2877 277 2899 283
rect 2964 277 3027 283
rect 3284 277 3315 283
rect 3482 276 3484 284
rect 3580 277 3604 283
rect 3796 277 3811 283
rect 4740 277 4771 283
rect 5476 277 5491 283
rect 5556 277 5571 283
rect 5620 277 5635 283
rect 5773 277 5788 283
rect 6317 277 6332 283
rect 285 257 323 263
rect 509 257 515 276
rect 2676 257 2691 263
rect 3124 257 3139 263
rect 4052 256 4060 264
rect 5309 257 5331 263
rect 5444 256 5452 264
rect 5668 257 5683 263
rect 628 236 630 244
rect 1620 236 1622 244
rect 2088 236 2092 244
rect 2938 214 2950 216
rect 5946 214 5958 216
rect 2923 206 2925 214
rect 2933 206 2935 214
rect 2943 206 2945 214
rect 2953 206 2955 214
rect 2963 206 2965 214
rect 5931 206 5933 214
rect 5941 206 5943 214
rect 5951 206 5953 214
rect 5961 206 5963 214
rect 5971 206 5973 214
rect 2938 204 2950 206
rect 5946 204 5958 206
rect 196 176 198 184
rect 1172 176 1176 184
rect 1268 176 1270 184
rect 1338 176 1340 184
rect 1652 176 1656 184
rect 2026 176 2028 184
rect 2458 176 2460 184
rect 4724 176 4726 184
rect 4820 176 4822 184
rect 1725 157 1740 163
rect 2909 157 2972 163
rect 3988 156 3996 164
rect 6045 157 6083 163
rect 157 143 163 156
rect 157 137 179 143
rect 269 137 284 143
rect 413 143 419 156
rect 397 137 419 143
rect 1117 137 1132 143
rect 1357 137 1436 143
rect 1917 137 1955 143
rect 2061 137 2099 143
rect 2324 137 2339 143
rect 2797 137 2835 143
rect 132 117 147 123
rect 637 117 659 123
rect 637 104 643 117
rect 781 117 819 123
rect 845 117 860 123
rect 925 117 963 123
rect 1080 117 1116 123
rect 1565 117 1587 123
rect 2045 117 2067 123
rect 2148 117 2179 123
rect 2381 117 2435 123
rect 2589 123 2595 136
rect 2797 124 2803 137
rect 3420 137 3444 143
rect 4093 137 4147 143
rect 4541 137 4556 143
rect 5076 137 5091 143
rect 5124 137 5139 143
rect 5284 137 5300 143
rect 6100 137 6116 143
rect 2573 117 2595 123
rect 2692 117 2707 123
rect 2749 117 2764 123
rect 2877 117 2899 123
rect 2916 117 2995 123
rect 3837 117 3852 123
rect 4061 117 4076 123
rect 4429 117 4492 123
rect 5588 117 5603 123
rect 6365 117 6396 123
rect 125 97 147 103
rect 324 97 339 103
rect 589 97 604 103
rect 813 97 835 103
rect 973 97 995 103
rect 1293 97 1331 103
rect 2429 97 2451 103
rect 4781 97 4796 103
rect 381 77 396 83
rect 1476 76 1480 84
rect 2269 77 2284 83
rect 1434 14 1446 16
rect 4442 14 4454 16
rect 1419 6 1421 14
rect 1429 6 1431 14
rect 1439 6 1441 14
rect 1449 6 1451 14
rect 1459 6 1461 14
rect 4427 6 4429 14
rect 4437 6 4439 14
rect 4447 6 4449 14
rect 4457 6 4459 14
rect 4467 6 4469 14
rect 1434 4 1446 6
rect 4442 4 4454 6
<< m2contact >>
rect 2915 5406 2923 5414
rect 2925 5406 2933 5414
rect 2935 5406 2943 5414
rect 2945 5406 2953 5414
rect 2955 5406 2963 5414
rect 2965 5406 2973 5414
rect 5923 5406 5931 5414
rect 5933 5406 5941 5414
rect 5943 5406 5951 5414
rect 5953 5406 5961 5414
rect 5963 5406 5971 5414
rect 5973 5406 5981 5414
rect 508 5376 516 5384
rect 604 5376 612 5384
rect 1100 5376 1108 5384
rect 1260 5376 1268 5384
rect 1548 5376 1556 5384
rect 2284 5376 2292 5384
rect 2572 5376 2580 5384
rect 2588 5376 2596 5384
rect 2812 5376 2820 5384
rect 2860 5376 2868 5384
rect 3612 5376 3620 5384
rect 3660 5376 3668 5384
rect 3708 5376 3716 5384
rect 3724 5376 3732 5384
rect 4204 5376 4212 5384
rect 4700 5376 4708 5384
rect 5436 5376 5444 5384
rect 5996 5376 6004 5384
rect 6604 5376 6612 5384
rect 6796 5376 6804 5384
rect 7052 5376 7060 5384
rect 7212 5376 7220 5384
rect 252 5356 260 5364
rect 492 5356 500 5364
rect 524 5356 532 5364
rect 540 5356 548 5364
rect 620 5356 628 5364
rect 796 5356 804 5364
rect 812 5356 820 5364
rect 844 5356 852 5364
rect 284 5336 292 5344
rect 316 5336 324 5344
rect 380 5336 388 5344
rect 396 5336 404 5344
rect 428 5336 436 5344
rect 668 5336 676 5344
rect 764 5336 772 5344
rect 796 5336 804 5344
rect 892 5356 900 5364
rect 1212 5356 1220 5364
rect 1276 5356 1284 5364
rect 1404 5356 1412 5364
rect 1484 5356 1492 5364
rect 1612 5356 1620 5364
rect 1836 5356 1844 5364
rect 1900 5356 1908 5364
rect 1996 5356 2004 5364
rect 2012 5356 2020 5364
rect 2332 5356 2340 5364
rect 3404 5356 3412 5364
rect 3916 5356 3924 5364
rect 4588 5356 4596 5364
rect 5676 5356 5684 5364
rect 6188 5356 6196 5364
rect 6988 5356 6996 5364
rect 908 5336 916 5344
rect 956 5336 964 5344
rect 1020 5336 1028 5344
rect 1084 5336 1092 5344
rect 1324 5336 1332 5344
rect 1356 5336 1364 5344
rect 1564 5336 1572 5344
rect 1596 5336 1604 5344
rect 1628 5336 1636 5344
rect 1644 5336 1652 5344
rect 1708 5336 1716 5344
rect 1756 5336 1764 5344
rect 1932 5336 1940 5344
rect 1964 5336 1972 5344
rect 2028 5336 2036 5344
rect 2092 5336 2100 5344
rect 2108 5336 2116 5344
rect 2204 5336 2212 5344
rect 2220 5336 2228 5344
rect 2316 5336 2324 5344
rect 2380 5336 2388 5344
rect 2748 5336 2756 5344
rect 3100 5336 3108 5344
rect 3324 5336 3332 5344
rect 3420 5336 3428 5344
rect 3452 5336 3460 5344
rect 3548 5336 3556 5344
rect 3884 5336 3892 5344
rect 3948 5336 3956 5344
rect 3996 5336 4004 5344
rect 4092 5336 4100 5344
rect 4220 5336 4228 5344
rect 4316 5336 4324 5344
rect 4652 5336 4660 5344
rect 4668 5336 4676 5344
rect 4812 5336 4820 5344
rect 4988 5336 4996 5344
rect 5052 5336 5060 5344
rect 5084 5336 5092 5344
rect 5260 5336 5268 5344
rect 5292 5336 5300 5344
rect 5356 5336 5364 5344
rect 5596 5336 5604 5344
rect 5628 5336 5636 5344
rect 5724 5336 5732 5344
rect 6060 5336 6068 5344
rect 6156 5336 6164 5344
rect 6220 5336 6228 5344
rect 6268 5336 6276 5344
rect 6492 5336 6500 5344
rect 6588 5336 6596 5344
rect 6764 5336 6772 5344
rect 6956 5336 6964 5344
rect 7068 5336 7076 5344
rect 44 5316 52 5324
rect 108 5316 116 5324
rect 204 5316 212 5324
rect 316 5316 324 5324
rect 380 5316 388 5324
rect 460 5316 468 5324
rect 572 5316 580 5324
rect 652 5316 660 5324
rect 700 5296 708 5304
rect 748 5316 756 5324
rect 764 5316 772 5324
rect 844 5316 852 5324
rect 972 5316 980 5324
rect 988 5316 996 5324
rect 1036 5316 1044 5324
rect 1052 5316 1060 5324
rect 1068 5316 1076 5324
rect 1164 5316 1172 5324
rect 1180 5316 1188 5324
rect 1228 5316 1236 5324
rect 1516 5316 1524 5324
rect 1660 5316 1668 5324
rect 1692 5316 1700 5324
rect 1004 5296 1012 5304
rect 1500 5296 1508 5304
rect 1596 5296 1604 5304
rect 1788 5316 1796 5324
rect 1852 5316 1860 5324
rect 1868 5316 1876 5324
rect 1916 5316 1924 5324
rect 2044 5316 2052 5324
rect 2076 5316 2084 5324
rect 2092 5316 2100 5324
rect 2140 5316 2148 5324
rect 2172 5316 2180 5324
rect 2364 5316 2372 5324
rect 2428 5316 2436 5324
rect 2524 5316 2532 5324
rect 2540 5316 2548 5324
rect 2716 5318 2724 5326
rect 2780 5316 2788 5324
rect 2828 5316 2836 5324
rect 3068 5318 3076 5326
rect 3212 5316 3220 5324
rect 3260 5318 3268 5326
rect 3340 5316 3348 5324
rect 3452 5316 3460 5324
rect 3468 5316 3476 5324
rect 3500 5316 3508 5324
rect 3564 5316 3572 5324
rect 3580 5316 3588 5324
rect 3628 5316 3636 5324
rect 3676 5316 3684 5324
rect 3852 5318 3860 5326
rect 3948 5316 3956 5324
rect 4012 5316 4020 5324
rect 4108 5316 4116 5324
rect 4236 5316 4244 5324
rect 4252 5316 4260 5324
rect 1932 5296 1940 5304
rect 2156 5296 2164 5304
rect 3372 5296 3380 5304
rect 3500 5296 3508 5304
rect 4348 5316 4356 5324
rect 4396 5316 4404 5324
rect 4492 5316 4500 5324
rect 4508 5316 4516 5324
rect 4556 5316 4564 5324
rect 4572 5316 4580 5324
rect 4620 5316 4628 5324
rect 4684 5316 4692 5324
rect 4796 5316 4804 5324
rect 4908 5316 4916 5324
rect 4956 5316 4964 5324
rect 4972 5316 4980 5324
rect 5004 5316 5012 5324
rect 4284 5296 4292 5304
rect 4924 5296 4932 5304
rect 5196 5316 5204 5324
rect 5308 5316 5316 5324
rect 5340 5316 5348 5324
rect 5388 5316 5396 5324
rect 5404 5316 5412 5324
rect 5516 5316 5524 5324
rect 5564 5318 5572 5326
rect 5052 5296 5060 5304
rect 5308 5296 5316 5304
rect 5372 5296 5380 5304
rect 5660 5296 5668 5304
rect 5708 5316 5716 5324
rect 5756 5316 5764 5324
rect 5804 5316 5812 5324
rect 5820 5316 5828 5324
rect 5852 5316 5860 5324
rect 5900 5316 5908 5324
rect 5916 5316 5924 5324
rect 6124 5318 6132 5326
rect 6220 5316 6228 5324
rect 6284 5316 6292 5324
rect 6316 5316 6324 5324
rect 6364 5316 6372 5324
rect 6380 5316 6388 5324
rect 6412 5316 6420 5324
rect 6460 5316 6468 5324
rect 6476 5316 6484 5324
rect 5772 5296 5780 5304
rect 6524 5296 6532 5304
rect 6572 5316 6580 5324
rect 6716 5316 6724 5324
rect 6924 5318 6932 5326
rect 7164 5336 7172 5344
rect 7196 5336 7204 5344
rect 7020 5316 7028 5324
rect 7084 5316 7092 5324
rect 7100 5316 7108 5324
rect 7276 5316 7284 5324
rect 7308 5316 7316 5324
rect 7164 5296 7172 5304
rect 12 5276 20 5284
rect 1484 5276 1492 5284
rect 1804 5276 1812 5284
rect 2940 5276 2948 5284
rect 5084 5276 5092 5284
rect 6572 5276 6580 5284
rect 748 5256 756 5264
rect 1132 5256 1140 5264
rect 1692 5256 1700 5264
rect 6428 5256 6436 5264
rect 60 5236 68 5244
rect 140 5236 148 5244
rect 156 5236 164 5244
rect 236 5236 244 5244
rect 300 5236 308 5244
rect 396 5236 404 5244
rect 460 5236 468 5244
rect 556 5236 564 5244
rect 860 5236 868 5244
rect 940 5236 948 5244
rect 1324 5236 1332 5244
rect 1820 5236 1828 5244
rect 2060 5236 2068 5244
rect 2364 5236 2372 5244
rect 2492 5236 2500 5244
rect 3132 5236 3140 5244
rect 4380 5236 4388 5244
rect 4540 5236 4548 5244
rect 5868 5236 5876 5244
rect 6332 5236 6340 5244
rect 1411 5206 1419 5214
rect 1421 5206 1429 5214
rect 1431 5206 1439 5214
rect 1441 5206 1449 5214
rect 1451 5206 1459 5214
rect 1461 5206 1469 5214
rect 4419 5206 4427 5214
rect 4429 5206 4437 5214
rect 4439 5206 4447 5214
rect 4449 5206 4457 5214
rect 4459 5206 4467 5214
rect 4469 5206 4477 5214
rect 1820 5176 1828 5184
rect 2268 5176 2276 5184
rect 2524 5176 2532 5184
rect 2540 5176 2548 5184
rect 3004 5176 3012 5184
rect 3804 5176 3812 5184
rect 5020 5176 5028 5184
rect 5372 5176 5380 5184
rect 6124 5176 6132 5184
rect 1100 5156 1108 5164
rect 348 5136 356 5144
rect 412 5136 420 5144
rect 2924 5136 2932 5144
rect 3052 5136 3060 5144
rect 3244 5136 3252 5144
rect 3596 5136 3604 5144
rect 3884 5136 3892 5144
rect 5308 5136 5316 5144
rect 5772 5136 5780 5144
rect 5884 5136 5892 5144
rect 6300 5136 6308 5144
rect 6332 5136 6340 5144
rect 6636 5136 6644 5144
rect 6828 5136 6836 5144
rect 6988 5136 6996 5144
rect 300 5116 308 5124
rect 380 5116 388 5124
rect 604 5116 612 5124
rect 636 5116 644 5124
rect 988 5116 996 5124
rect 1052 5116 1060 5124
rect 1148 5116 1156 5124
rect 1164 5116 1172 5124
rect 1868 5116 1876 5124
rect 1932 5116 1940 5124
rect 2156 5116 2164 5124
rect 2172 5116 2180 5124
rect 2348 5116 2356 5124
rect 2460 5116 2468 5124
rect 2780 5116 2788 5124
rect 3484 5116 3492 5124
rect 140 5096 148 5104
rect 188 5096 196 5104
rect 300 5096 308 5104
rect 332 5096 340 5104
rect 396 5096 404 5104
rect 460 5096 468 5104
rect 492 5096 500 5104
rect 524 5096 532 5104
rect 556 5096 564 5104
rect 588 5096 596 5104
rect 684 5096 692 5104
rect 748 5096 756 5104
rect 796 5096 804 5104
rect 876 5096 884 5104
rect 924 5096 932 5104
rect 940 5096 948 5104
rect 1020 5096 1028 5104
rect 1036 5096 1044 5104
rect 1100 5096 1108 5104
rect 1148 5096 1156 5104
rect 1212 5096 1220 5104
rect 1228 5096 1236 5104
rect 1260 5096 1268 5104
rect 1308 5096 1316 5104
rect 1372 5096 1380 5104
rect 1484 5096 1492 5104
rect 1548 5096 1556 5104
rect 1596 5096 1604 5104
rect 1644 5096 1652 5104
rect 1772 5096 1780 5104
rect 1836 5096 1844 5104
rect 1900 5096 1908 5104
rect 2060 5096 2068 5104
rect 2108 5096 2116 5104
rect 2156 5096 2164 5104
rect 2204 5096 2212 5104
rect 2236 5096 2244 5104
rect 2284 5096 2292 5104
rect 2428 5096 2436 5104
rect 2476 5096 2484 5104
rect 2716 5094 2724 5102
rect 2828 5096 2836 5104
rect 2860 5096 2868 5104
rect 2892 5096 2900 5104
rect 3036 5096 3044 5104
rect 3116 5096 3124 5104
rect 3148 5096 3156 5104
rect 3308 5096 3316 5104
rect 3372 5094 3380 5102
rect 3452 5096 3460 5104
rect 3484 5096 3492 5104
rect 3548 5096 3556 5104
rect 3564 5096 3572 5104
rect 3740 5094 3748 5102
rect 3836 5096 3844 5104
rect 3980 5094 3988 5102
rect 4108 5096 4116 5104
rect 4252 5096 4260 5104
rect 4268 5096 4276 5104
rect 4300 5116 4308 5124
rect 4652 5116 4660 5124
rect 4460 5094 4468 5102
rect 4620 5096 4628 5104
rect 4684 5096 4692 5104
rect 4700 5096 4708 5104
rect 4748 5096 4756 5104
rect 4764 5096 4772 5104
rect 4796 5096 4804 5104
rect 4860 5096 4868 5104
rect 4892 5096 4900 5104
rect 4956 5096 4964 5104
rect 5052 5096 5060 5104
rect 5164 5116 5172 5124
rect 5244 5116 5252 5124
rect 5436 5116 5444 5124
rect 5116 5096 5124 5104
rect 5148 5096 5156 5104
rect 5212 5096 5220 5104
rect 5244 5096 5252 5104
rect 5308 5096 5316 5104
rect 5356 5096 5364 5104
rect 5404 5096 5412 5104
rect 5420 5096 5428 5104
rect 5468 5096 5476 5104
rect 5500 5096 5508 5104
rect 5932 5116 5940 5124
rect 7228 5116 7236 5124
rect 7356 5116 7364 5124
rect 5580 5096 5588 5104
rect 5692 5096 5700 5104
rect 5772 5096 5780 5104
rect 5788 5096 5796 5104
rect 5836 5096 5844 5104
rect 5884 5096 5892 5104
rect 5996 5096 6004 5104
rect 6012 5096 6020 5104
rect 6108 5096 6116 5104
rect 6156 5096 6164 5104
rect 6172 5096 6180 5104
rect 6188 5096 6196 5104
rect 6284 5096 6292 5104
rect 6412 5096 6420 5104
rect 6524 5096 6532 5104
rect 6556 5096 6564 5104
rect 6588 5096 6596 5104
rect 6716 5096 6724 5104
rect 6908 5096 6916 5104
rect 7116 5094 7124 5102
rect 7212 5096 7220 5104
rect 7276 5096 7284 5104
rect 7308 5096 7316 5104
rect 12 5076 20 5084
rect 108 5076 116 5084
rect 124 5076 132 5084
rect 300 5076 308 5084
rect 444 5076 452 5084
rect 508 5076 516 5084
rect 540 5076 548 5084
rect 604 5076 612 5084
rect 636 5076 644 5084
rect 716 5076 724 5084
rect 732 5076 740 5084
rect 828 5076 836 5084
rect 940 5076 948 5084
rect 1004 5076 1012 5084
rect 1116 5076 1124 5084
rect 1148 5076 1156 5084
rect 1212 5076 1220 5084
rect 1356 5076 1364 5084
rect 1500 5076 1508 5084
rect 1692 5076 1700 5084
rect 1724 5076 1732 5084
rect 1788 5076 1796 5084
rect 1884 5076 1892 5084
rect 1916 5076 1924 5084
rect 1964 5076 1972 5084
rect 2044 5076 2052 5084
rect 2108 5076 2116 5084
rect 2220 5076 2228 5084
rect 2300 5076 2308 5084
rect 2380 5076 2388 5084
rect 2412 5076 2420 5084
rect 2444 5076 2452 5084
rect 2748 5076 2756 5084
rect 2812 5076 2820 5084
rect 2876 5076 2884 5084
rect 3212 5076 3220 5084
rect 3436 5076 3444 5084
rect 3532 5076 3540 5084
rect 3772 5076 3780 5084
rect 4236 5076 4244 5084
rect 4332 5076 4340 5084
rect 4492 5076 4500 5084
rect 4604 5076 4612 5084
rect 4668 5076 4676 5084
rect 4780 5076 4788 5084
rect 4844 5076 4852 5084
rect 4892 5076 4900 5084
rect 5004 5076 5012 5084
rect 5068 5076 5076 5084
rect 5084 5076 5092 5084
rect 5132 5076 5140 5084
rect 5196 5076 5204 5084
rect 5324 5076 5332 5084
rect 5484 5076 5492 5084
rect 5548 5076 5556 5084
rect 5564 5076 5572 5084
rect 5596 5076 5604 5084
rect 5628 5076 5636 5084
rect 5788 5076 5796 5084
rect 5820 5076 5828 5084
rect 5852 5076 5860 5084
rect 5868 5076 5876 5084
rect 220 5056 228 5064
rect 236 5056 244 5064
rect 428 5056 436 5064
rect 668 5056 676 5064
rect 828 5056 836 5064
rect 1068 5056 1076 5064
rect 1260 5056 1268 5064
rect 1292 5056 1300 5064
rect 1340 5056 1348 5064
rect 1596 5056 1604 5064
rect 1628 5056 1636 5064
rect 1692 5056 1700 5064
rect 1804 5056 1812 5064
rect 1852 5056 1860 5064
rect 1980 5056 1988 5064
rect 2092 5056 2100 5064
rect 2332 5056 2340 5064
rect 2364 5056 2372 5064
rect 2476 5056 2484 5064
rect 2540 5056 2548 5064
rect 3740 5056 3748 5064
rect 4092 5056 4100 5064
rect 4860 5056 4868 5064
rect 4908 5056 4916 5064
rect 4988 5056 4996 5064
rect 5180 5056 5188 5064
rect 5644 5056 5652 5064
rect 5724 5056 5732 5064
rect 6028 5056 6036 5064
rect 6220 5056 6228 5064
rect 6268 5076 6276 5084
rect 6460 5076 6468 5084
rect 6572 5076 6580 5084
rect 6764 5076 6772 5084
rect 6956 5076 6964 5084
rect 7148 5076 7156 5084
rect 7260 5076 7268 5084
rect 7292 5076 7300 5084
rect 6252 5056 6260 5064
rect 6492 5056 6500 5064
rect 7180 5056 7188 5064
rect 60 5036 68 5044
rect 172 5036 180 5044
rect 204 5036 212 5044
rect 364 5036 372 5044
rect 492 5036 500 5044
rect 604 5036 612 5044
rect 780 5036 788 5044
rect 812 5036 820 5044
rect 892 5036 900 5044
rect 988 5036 996 5044
rect 1244 5036 1252 5044
rect 1404 5036 1412 5044
rect 1516 5036 1524 5044
rect 1612 5036 1620 5044
rect 1772 5036 1780 5044
rect 1948 5036 1956 5044
rect 2028 5036 2036 5044
rect 2076 5036 2084 5044
rect 2156 5036 2164 5044
rect 2316 5036 2324 5044
rect 2588 5036 2596 5044
rect 3612 5036 3620 5044
rect 3852 5036 3860 5044
rect 4220 5036 4228 5044
rect 4588 5036 4596 5044
rect 4716 5036 4724 5044
rect 4796 5036 4804 5044
rect 4876 5036 4884 5044
rect 5436 5036 5444 5044
rect 5708 5036 5716 5044
rect 6604 5036 6612 5044
rect 6796 5036 6804 5044
rect 7340 5036 7348 5044
rect 2915 5006 2923 5014
rect 2925 5006 2933 5014
rect 2935 5006 2943 5014
rect 2945 5006 2953 5014
rect 2955 5006 2963 5014
rect 2965 5006 2973 5014
rect 5923 5006 5931 5014
rect 5933 5006 5941 5014
rect 5943 5006 5951 5014
rect 5953 5006 5961 5014
rect 5963 5006 5971 5014
rect 5973 5006 5981 5014
rect 76 4976 84 4984
rect 972 4976 980 4984
rect 1004 4976 1012 4984
rect 1484 4976 1492 4984
rect 1756 4976 1764 4984
rect 2236 4976 2244 4984
rect 2540 4976 2548 4984
rect 2636 4976 2644 4984
rect 2988 4976 2996 4984
rect 3388 4976 3396 4984
rect 3436 4976 3444 4984
rect 3532 4976 3540 4984
rect 3980 4976 3988 4984
rect 4044 4976 4052 4984
rect 4252 4976 4260 4984
rect 4284 4976 4292 4984
rect 4364 4976 4372 4984
rect 4668 4976 4676 4984
rect 4732 4976 4740 4984
rect 5020 4976 5028 4984
rect 5420 4976 5428 4984
rect 5676 4976 5684 4984
rect 6396 4976 6404 4984
rect 6636 4976 6644 4984
rect 7180 4976 7188 4984
rect 204 4956 212 4964
rect 252 4956 260 4964
rect 540 4956 548 4964
rect 684 4956 692 4964
rect 716 4956 724 4964
rect 812 4956 820 4964
rect 876 4956 884 4964
rect 908 4956 916 4964
rect 1132 4956 1140 4964
rect 1196 4956 1204 4964
rect 1228 4956 1236 4964
rect 1516 4956 1524 4964
rect 1532 4956 1540 4964
rect 1660 4956 1668 4964
rect 1676 4956 1684 4964
rect 1804 4956 1812 4964
rect 1996 4956 2004 4964
rect 2076 4956 2084 4964
rect 2220 4956 2228 4964
rect 2252 4956 2260 4964
rect 2300 4956 2308 4964
rect 2316 4956 2324 4964
rect 2380 4956 2388 4964
rect 2412 4956 2420 4964
rect 2604 4956 2612 4964
rect 2684 4956 2692 4964
rect 2732 4956 2740 4964
rect 2828 4956 2836 4964
rect 3964 4956 3972 4964
rect 4268 4956 4276 4964
rect 4428 4956 4436 4964
rect 4556 4956 4564 4964
rect 5068 4956 5076 4964
rect 12 4936 20 4944
rect 124 4936 132 4944
rect 252 4936 260 4944
rect 316 4936 324 4944
rect 572 4936 580 4944
rect 588 4936 596 4944
rect 604 4936 612 4944
rect 668 4936 676 4944
rect 812 4936 820 4944
rect 940 4936 948 4944
rect 988 4936 996 4944
rect 1052 4936 1060 4944
rect 1068 4936 1076 4944
rect 1164 4936 1172 4944
rect 1196 4936 1204 4944
rect 1228 4936 1236 4944
rect 1292 4936 1300 4944
rect 1372 4936 1380 4944
rect 1580 4936 1588 4944
rect 1612 4936 1620 4944
rect 1708 4936 1716 4944
rect 1820 4936 1828 4944
rect 1884 4936 1892 4944
rect 1900 4936 1908 4944
rect 1996 4936 2004 4944
rect 2108 4936 2116 4944
rect 2188 4936 2196 4944
rect 2460 4936 2468 4944
rect 2524 4936 2532 4944
rect 2572 4936 2580 4944
rect 2588 4936 2596 4944
rect 2620 4936 2628 4944
rect 2892 4936 2900 4944
rect 3052 4936 3060 4944
rect 3100 4936 3108 4944
rect 3132 4936 3140 4944
rect 3180 4936 3188 4944
rect 3276 4936 3284 4944
rect 3292 4936 3300 4944
rect 3404 4936 3412 4944
rect 3580 4936 3588 4944
rect 3676 4936 3684 4944
rect 3916 4936 3924 4944
rect 3948 4936 3956 4944
rect 3996 4936 4004 4944
rect 4060 4936 4068 4944
rect 4092 4936 4100 4944
rect 4300 4936 4308 4944
rect 4348 4936 4356 4944
rect 4444 4936 4452 4944
rect 4604 4936 4612 4944
rect 4620 4936 4628 4944
rect 4684 4936 4692 4944
rect 4764 4936 4772 4944
rect 4860 4936 4868 4944
rect 5692 4956 5700 4964
rect 6012 4956 6020 4964
rect 6140 4956 6148 4964
rect 6556 4956 6564 4964
rect 6588 4956 6596 4964
rect 6652 4956 6660 4964
rect 6908 4956 6916 4964
rect 6940 4956 6948 4964
rect 5116 4936 5124 4944
rect 5164 4936 5172 4944
rect 5436 4936 5444 4944
rect 5516 4936 5524 4944
rect 5724 4936 5732 4944
rect 5740 4936 5748 4944
rect 5804 4936 5812 4944
rect 6028 4936 6036 4944
rect 6092 4936 6100 4944
rect 6156 4936 6164 4944
rect 6188 4936 6196 4944
rect 6220 4936 6228 4944
rect 6284 4936 6292 4944
rect 6348 4936 6356 4944
rect 6460 4936 6468 4944
rect 108 4916 116 4924
rect 140 4916 148 4924
rect 156 4916 164 4924
rect 220 4916 228 4924
rect 300 4916 308 4924
rect 348 4916 356 4924
rect 396 4916 404 4924
rect 412 4916 420 4924
rect 492 4916 500 4924
rect 620 4916 628 4924
rect 764 4916 772 4924
rect 780 4916 788 4924
rect 860 4916 868 4924
rect 940 4916 948 4924
rect 1004 4916 1012 4924
rect 1036 4916 1044 4924
rect 1100 4916 1108 4924
rect 1116 4916 1124 4924
rect 1148 4916 1156 4924
rect 1276 4916 1284 4924
rect 1324 4916 1332 4924
rect 1436 4916 1444 4924
rect 1596 4916 1604 4924
rect 1756 4916 1764 4924
rect 1836 4916 1844 4924
rect 1868 4916 1876 4924
rect 1916 4916 1924 4924
rect 2044 4916 2052 4924
rect 2092 4916 2100 4924
rect 2124 4916 2132 4924
rect 2156 4916 2164 4924
rect 2172 4916 2180 4924
rect 2268 4916 2276 4924
rect 2364 4916 2372 4924
rect 2412 4916 2420 4924
rect 2460 4916 2468 4924
rect 2476 4916 2484 4924
rect 2508 4916 2516 4924
rect 172 4896 180 4904
rect 508 4896 516 4904
rect 972 4896 980 4904
rect 1244 4896 1252 4904
rect 1308 4896 1316 4904
rect 1372 4896 1380 4904
rect 1948 4896 1956 4904
rect 2044 4896 2052 4904
rect 2156 4896 2164 4904
rect 2476 4896 2484 4904
rect 2700 4916 2708 4924
rect 2780 4916 2788 4924
rect 2796 4916 2804 4924
rect 2844 4916 2852 4924
rect 2924 4896 2932 4904
rect 3036 4916 3044 4924
rect 3084 4916 3092 4924
rect 3196 4916 3204 4924
rect 3308 4916 3316 4924
rect 3324 4916 3332 4924
rect 3420 4916 3428 4924
rect 3468 4916 3476 4924
rect 3516 4916 3524 4924
rect 3564 4916 3572 4924
rect 3580 4916 3588 4924
rect 3660 4916 3668 4924
rect 3692 4916 3700 4924
rect 3772 4916 3780 4924
rect 3820 4916 3828 4924
rect 3932 4916 3940 4924
rect 4012 4916 4020 4924
rect 4140 4916 4148 4924
rect 4188 4916 4196 4924
rect 4316 4916 4324 4924
rect 4332 4916 4340 4924
rect 4396 4916 4404 4924
rect 3164 4896 3172 4904
rect 3228 4896 3236 4904
rect 3244 4896 3252 4904
rect 3356 4896 3364 4904
rect 3628 4896 3636 4904
rect 3900 4896 3908 4904
rect 4540 4896 4548 4904
rect 4604 4916 4612 4924
rect 4620 4916 4628 4924
rect 4684 4916 4692 4924
rect 4748 4916 4756 4924
rect 4812 4916 4820 4924
rect 4828 4916 4836 4924
rect 4908 4916 4916 4924
rect 5036 4916 5044 4924
rect 5068 4916 5076 4924
rect 5132 4916 5140 4924
rect 5164 4916 5172 4924
rect 5212 4916 5220 4924
rect 5228 4916 5236 4924
rect 5308 4916 5316 4924
rect 5356 4916 5364 4924
rect 5452 4916 5460 4924
rect 5468 4916 5476 4924
rect 5580 4916 5588 4924
rect 5740 4916 5748 4924
rect 5756 4916 5764 4924
rect 5788 4916 5796 4924
rect 5820 4916 5828 4924
rect 5836 4916 5844 4924
rect 5884 4916 5892 4924
rect 5964 4916 5972 4924
rect 6076 4916 6084 4924
rect 6108 4916 6116 4924
rect 6204 4916 6212 4924
rect 4668 4896 4676 4904
rect 4732 4896 4740 4904
rect 5484 4896 5492 4904
rect 5788 4896 5796 4904
rect 6268 4916 6276 4924
rect 6300 4916 6308 4924
rect 6332 4916 6340 4924
rect 6380 4916 6388 4924
rect 6428 4916 6436 4924
rect 6444 4916 6452 4924
rect 6476 4916 6484 4924
rect 6524 4916 6532 4924
rect 6540 4916 6548 4924
rect 6620 4936 6628 4944
rect 7052 4956 7060 4964
rect 6604 4916 6612 4924
rect 6668 4916 6676 4924
rect 6684 4916 6692 4924
rect 6732 4916 6740 4924
rect 6764 4916 6772 4924
rect 6780 4916 6788 4924
rect 6828 4916 6836 4924
rect 6860 4916 6868 4924
rect 6988 4936 6996 4944
rect 6972 4916 6980 4924
rect 7004 4916 7012 4924
rect 7100 4936 7108 4944
rect 7164 4936 7172 4944
rect 7116 4916 7124 4924
rect 7244 4916 7252 4924
rect 7292 4916 7300 4924
rect 6300 4896 6308 4904
rect 7132 4896 7140 4904
rect 476 4876 484 4884
rect 636 4876 644 4884
rect 1340 4876 1348 4884
rect 2028 4876 2036 4884
rect 2428 4876 2436 4884
rect 2892 4876 2900 4884
rect 3484 4876 3492 4884
rect 5868 4876 5876 4884
rect 6268 4876 6276 4884
rect 1324 4856 1332 4864
rect 2316 4856 2324 4864
rect 188 4836 196 4844
rect 236 4836 244 4844
rect 364 4836 372 4844
rect 428 4836 436 4844
rect 732 4836 740 4844
rect 796 4836 804 4844
rect 892 4836 900 4844
rect 1196 4836 1204 4844
rect 1868 4836 1876 4844
rect 1980 4836 1988 4844
rect 2044 4836 2052 4844
rect 2204 4836 2212 4844
rect 2300 4836 2308 4844
rect 2732 4836 2740 4844
rect 2748 4836 2756 4844
rect 3708 4836 3716 4844
rect 5676 4836 5684 4844
rect 6044 4836 6052 4844
rect 6700 4836 6708 4844
rect 6796 4836 6804 4844
rect 7068 4836 7076 4844
rect 7148 4836 7156 4844
rect 1411 4806 1419 4814
rect 1421 4806 1429 4814
rect 1431 4806 1439 4814
rect 1441 4806 1449 4814
rect 1451 4806 1459 4814
rect 1461 4806 1469 4814
rect 4419 4806 4427 4814
rect 4429 4806 4437 4814
rect 4439 4806 4447 4814
rect 4449 4806 4457 4814
rect 4459 4806 4467 4814
rect 4469 4806 4477 4814
rect 2604 4776 2612 4784
rect 3164 4776 3172 4784
rect 3420 4776 3428 4784
rect 3452 4776 3460 4784
rect 3468 4776 3476 4784
rect 3852 4776 3860 4784
rect 5260 4776 5268 4784
rect 5308 4776 5316 4784
rect 5788 4776 5796 4784
rect 5916 4776 5924 4784
rect 6268 4776 6276 4784
rect 6972 4776 6980 4784
rect 4620 4756 4628 4764
rect 5132 4756 5140 4764
rect 5868 4756 5876 4764
rect 6108 4756 6116 4764
rect 1116 4736 1124 4744
rect 2140 4736 2148 4744
rect 2204 4736 2212 4744
rect 2668 4736 2676 4744
rect 5212 4736 5220 4744
rect 5548 4736 5556 4744
rect 5660 4736 5668 4744
rect 6076 4736 6084 4744
rect 6588 4736 6596 4744
rect 188 4716 196 4724
rect 460 4716 468 4724
rect 476 4716 484 4724
rect 1052 4716 1060 4724
rect 1308 4716 1316 4724
rect 1468 4716 1476 4724
rect 44 4696 52 4704
rect 252 4696 260 4704
rect 284 4696 292 4704
rect 156 4676 164 4684
rect 332 4696 340 4704
rect 380 4696 388 4704
rect 428 4696 436 4704
rect 556 4696 564 4704
rect 620 4696 628 4704
rect 844 4696 852 4704
rect 876 4696 884 4704
rect 892 4696 900 4704
rect 988 4696 996 4704
rect 1004 4696 1012 4704
rect 1100 4696 1108 4704
rect 1260 4696 1268 4704
rect 1292 4696 1300 4704
rect 1356 4696 1364 4704
rect 1372 4696 1380 4704
rect 1516 4696 1524 4704
rect 1612 4696 1620 4704
rect 1724 4696 1732 4704
rect 1740 4696 1748 4704
rect 2108 4716 2116 4724
rect 2172 4716 2180 4724
rect 2428 4716 2436 4724
rect 2588 4716 2596 4724
rect 2700 4716 2708 4724
rect 4108 4716 4116 4724
rect 4236 4716 4244 4724
rect 4652 4716 4660 4724
rect 1948 4696 1956 4704
rect 2028 4696 2036 4704
rect 2060 4696 2068 4704
rect 2092 4696 2100 4704
rect 2124 4696 2132 4704
rect 2204 4696 2212 4704
rect 2220 4696 2228 4704
rect 2300 4696 2308 4704
rect 2316 4696 2324 4704
rect 2380 4696 2388 4704
rect 2396 4696 2404 4704
rect 2492 4696 2500 4704
rect 2540 4696 2548 4704
rect 2572 4696 2580 4704
rect 2636 4696 2644 4704
rect 2684 4696 2692 4704
rect 2764 4696 2772 4704
rect 2844 4696 2852 4704
rect 2876 4696 2884 4704
rect 3212 4696 3220 4704
rect 3260 4696 3268 4704
rect 3500 4696 3508 4704
rect 3564 4696 3572 4704
rect 3660 4696 3668 4704
rect 3804 4696 3812 4704
rect 3996 4694 4004 4702
rect 4076 4696 4084 4704
rect 4124 4696 4132 4704
rect 4172 4696 4180 4704
rect 4204 4696 4212 4704
rect 4268 4696 4276 4704
rect 4284 4696 4292 4704
rect 4364 4696 4372 4704
rect 4508 4696 4516 4704
rect 4636 4696 4644 4704
rect 4700 4716 4708 4724
rect 4956 4716 4964 4724
rect 4876 4694 4884 4702
rect 4956 4696 4964 4704
rect 5004 4716 5012 4724
rect 5084 4716 5092 4724
rect 5244 4716 5252 4724
rect 5036 4696 5044 4704
rect 5100 4696 5108 4704
rect 5132 4696 5140 4704
rect 5180 4696 5188 4704
rect 5212 4696 5220 4704
rect 5292 4696 5300 4704
rect 5340 4696 5348 4704
rect 5484 4694 5492 4702
rect 5564 4696 5572 4704
rect 5628 4696 5636 4704
rect 6172 4716 6180 4724
rect 6412 4716 6420 4724
rect 5692 4696 5700 4704
rect 5708 4696 5716 4704
rect 5772 4696 5780 4704
rect 5820 4696 5828 4704
rect 5836 4696 5844 4704
rect 5900 4696 5908 4704
rect 5948 4696 5956 4704
rect 5964 4696 5972 4704
rect 6076 4696 6084 4704
rect 6092 4696 6100 4704
rect 6140 4696 6148 4704
rect 6204 4696 6212 4704
rect 6252 4696 6260 4704
rect 6300 4696 6308 4704
rect 6316 4696 6324 4704
rect 6332 4696 6340 4704
rect 6364 4696 6372 4704
rect 6380 4696 6388 4704
rect 6428 4696 6436 4704
rect 6444 4696 6452 4704
rect 6508 4696 6516 4704
rect 6572 4696 6580 4704
rect 6700 4696 6708 4704
rect 6892 4696 6900 4704
rect 7084 4696 7092 4704
rect 7228 4696 7236 4704
rect 7276 4696 7284 4704
rect 364 4676 372 4684
rect 108 4656 116 4664
rect 140 4656 148 4664
rect 204 4656 212 4664
rect 236 4656 244 4664
rect 252 4656 260 4664
rect 284 4656 292 4664
rect 332 4656 340 4664
rect 364 4656 372 4664
rect 508 4676 516 4684
rect 572 4676 580 4684
rect 668 4676 676 4684
rect 796 4676 804 4684
rect 812 4676 820 4684
rect 892 4676 900 4684
rect 1004 4676 1012 4684
rect 460 4656 468 4664
rect 588 4656 596 4664
rect 620 4656 628 4664
rect 636 4656 644 4664
rect 716 4656 724 4664
rect 732 4656 740 4664
rect 812 4656 820 4664
rect 940 4656 948 4664
rect 956 4656 964 4664
rect 1100 4676 1108 4684
rect 1180 4656 1188 4664
rect 1244 4676 1252 4684
rect 1340 4676 1348 4684
rect 1516 4676 1524 4684
rect 1532 4676 1540 4684
rect 1628 4676 1636 4684
rect 1724 4676 1732 4684
rect 1756 4676 1764 4684
rect 1788 4676 1796 4684
rect 1836 4676 1844 4684
rect 1932 4676 1940 4684
rect 1996 4676 2004 4684
rect 2076 4676 2084 4684
rect 2332 4676 2340 4684
rect 2460 4676 2468 4684
rect 2540 4676 2548 4684
rect 2652 4676 2660 4684
rect 2828 4676 2836 4684
rect 1388 4656 1396 4664
rect 1564 4656 1572 4664
rect 1580 4656 1588 4664
rect 1772 4656 1780 4664
rect 1804 4656 1812 4664
rect 1996 4656 2004 4664
rect 2156 4656 2164 4664
rect 2252 4656 2260 4664
rect 2364 4656 2372 4664
rect 2412 4656 2420 4664
rect 2716 4656 2724 4664
rect 2780 4656 2788 4664
rect 2988 4676 2996 4684
rect 3004 4656 3012 4664
rect 3068 4676 3076 4684
rect 3276 4676 3284 4684
rect 3292 4676 3300 4684
rect 3388 4676 3396 4684
rect 3564 4676 3572 4684
rect 3692 4676 3700 4684
rect 3740 4676 3748 4684
rect 4028 4676 4036 4684
rect 4060 4676 4068 4684
rect 4156 4676 4164 4684
rect 4188 4676 4196 4684
rect 4300 4676 4308 4684
rect 4348 4676 4356 4684
rect 4636 4676 4644 4684
rect 4732 4676 4740 4684
rect 4844 4676 4852 4684
rect 4940 4676 4948 4684
rect 5052 4676 5060 4684
rect 5116 4676 5124 4684
rect 5180 4676 5188 4684
rect 5196 4676 5204 4684
rect 5516 4676 5524 4684
rect 5612 4676 5620 4684
rect 5724 4676 5732 4684
rect 6092 4676 6100 4684
rect 6156 4676 6164 4684
rect 6220 4676 6228 4684
rect 6332 4676 6340 4684
rect 6396 4676 6404 4684
rect 6476 4676 6484 4684
rect 6556 4676 6564 4684
rect 6748 4676 6756 4684
rect 6844 4676 6852 4684
rect 6940 4676 6948 4684
rect 7132 4676 7140 4684
rect 3132 4656 3140 4664
rect 3148 4656 3156 4664
rect 3180 4656 3188 4664
rect 3404 4656 3412 4664
rect 3436 4656 3444 4664
rect 3516 4656 3524 4664
rect 4236 4656 4244 4664
rect 4316 4656 4324 4664
rect 4492 4656 4500 4664
rect 4588 4656 4596 4664
rect 5068 4656 5076 4664
rect 5740 4656 5748 4664
rect 6028 4656 6036 4664
rect 6172 4656 6180 4664
rect 6540 4656 6548 4664
rect 12 4636 20 4644
rect 124 4636 132 4644
rect 188 4636 196 4644
rect 492 4636 500 4644
rect 524 4636 532 4644
rect 652 4636 660 4644
rect 748 4636 756 4644
rect 764 4636 772 4644
rect 924 4636 932 4644
rect 972 4636 980 4644
rect 1052 4636 1060 4644
rect 1068 4636 1076 4644
rect 1212 4636 1220 4644
rect 1292 4636 1300 4644
rect 1484 4636 1492 4644
rect 1548 4636 1556 4644
rect 2348 4636 2356 4644
rect 2428 4636 2436 4644
rect 2524 4636 2532 4644
rect 2732 4636 2740 4644
rect 3084 4636 3092 4644
rect 3228 4636 3236 4644
rect 3324 4636 3332 4644
rect 3532 4636 3540 4644
rect 3580 4636 3588 4644
rect 3772 4636 3780 4644
rect 3868 4636 3876 4644
rect 4332 4636 4340 4644
rect 4748 4636 4756 4644
rect 5308 4636 5316 4644
rect 5356 4636 5364 4644
rect 6780 4636 6788 4644
rect 7164 4636 7172 4644
rect 2915 4606 2923 4614
rect 2925 4606 2933 4614
rect 2935 4606 2943 4614
rect 2945 4606 2953 4614
rect 2955 4606 2963 4614
rect 2965 4606 2973 4614
rect 5923 4606 5931 4614
rect 5933 4606 5941 4614
rect 5943 4606 5951 4614
rect 5953 4606 5961 4614
rect 5963 4606 5971 4614
rect 5973 4606 5981 4614
rect 268 4576 276 4584
rect 1756 4576 1764 4584
rect 1852 4576 1860 4584
rect 1916 4576 1924 4584
rect 1964 4576 1972 4584
rect 2108 4576 2116 4584
rect 2604 4576 2612 4584
rect 2652 4576 2660 4584
rect 2684 4576 2692 4584
rect 3516 4576 3524 4584
rect 3548 4576 3556 4584
rect 3660 4576 3668 4584
rect 3708 4576 3716 4584
rect 3852 4576 3860 4584
rect 3964 4576 3972 4584
rect 4396 4576 4404 4584
rect 4540 4576 4548 4584
rect 4668 4576 4676 4584
rect 4732 4576 4740 4584
rect 4860 4576 4868 4584
rect 5260 4576 5268 4584
rect 5324 4576 5332 4584
rect 5532 4576 5540 4584
rect 5724 4576 5732 4584
rect 5772 4576 5780 4584
rect 5852 4576 5860 4584
rect 6012 4576 6020 4584
rect 6140 4576 6148 4584
rect 6236 4576 6244 4584
rect 6812 4576 6820 4584
rect 6924 4576 6932 4584
rect 7020 4576 7028 4584
rect 12 4556 20 4564
rect 76 4556 84 4564
rect 316 4556 324 4564
rect 396 4556 404 4564
rect 444 4556 452 4564
rect 620 4556 628 4564
rect 700 4556 708 4564
rect 764 4556 772 4564
rect 812 4556 820 4564
rect 828 4556 836 4564
rect 924 4556 932 4564
rect 972 4556 980 4564
rect 1036 4556 1044 4564
rect 1116 4556 1124 4564
rect 1132 4556 1140 4564
rect 1404 4556 1412 4564
rect 1596 4556 1604 4564
rect 1612 4556 1620 4564
rect 1868 4556 1876 4564
rect 2028 4556 2036 4564
rect 2060 4556 2068 4564
rect 2316 4556 2324 4564
rect 2412 4556 2420 4564
rect 2540 4556 2548 4564
rect 2620 4556 2628 4564
rect 2732 4556 2740 4564
rect 2860 4556 2868 4564
rect 3532 4556 3540 4564
rect 3644 4556 3652 4564
rect 3788 4556 3796 4564
rect 4508 4556 4516 4564
rect 140 4536 148 4544
rect 188 4536 196 4544
rect 44 4516 52 4524
rect 92 4516 100 4524
rect 124 4516 132 4524
rect 300 4536 308 4544
rect 348 4536 356 4544
rect 476 4536 484 4544
rect 684 4536 692 4544
rect 844 4536 852 4544
rect 1020 4536 1028 4544
rect 1084 4536 1092 4544
rect 1164 4536 1172 4544
rect 1180 4536 1188 4544
rect 1276 4536 1284 4544
rect 1324 4536 1332 4544
rect 1372 4532 1380 4540
rect 1388 4536 1396 4544
rect 1500 4536 1508 4544
rect 1564 4536 1572 4544
rect 1900 4536 1908 4544
rect 1932 4536 1940 4544
rect 2012 4536 2020 4544
rect 2060 4536 2068 4544
rect 2124 4536 2132 4544
rect 2140 4536 2148 4544
rect 2460 4536 2468 4544
rect 2540 4536 2548 4544
rect 2588 4536 2596 4544
rect 2668 4536 2676 4544
rect 2780 4536 2788 4544
rect 3020 4536 3028 4544
rect 3116 4536 3124 4544
rect 3132 4536 3140 4544
rect 3292 4536 3300 4544
rect 3388 4536 3396 4544
rect 3468 4536 3476 4544
rect 3564 4536 3572 4544
rect 3644 4536 3652 4544
rect 3676 4536 3684 4544
rect 3756 4536 3764 4544
rect 3804 4536 3812 4544
rect 3900 4536 3908 4544
rect 3980 4536 3988 4544
rect 4092 4536 4100 4544
rect 4188 4536 4196 4544
rect 4780 4556 4788 4564
rect 5468 4556 5476 4564
rect 5676 4556 5684 4564
rect 6028 4556 6036 4564
rect 6060 4556 6068 4564
rect 6108 4556 6116 4564
rect 6252 4556 6260 4564
rect 6748 4556 6756 4564
rect 6860 4556 6868 4564
rect 4556 4536 4564 4544
rect 4588 4536 4596 4544
rect 4636 4536 4644 4544
rect 4652 4536 4660 4544
rect 4716 4536 4724 4544
rect 4924 4536 4932 4544
rect 4956 4536 4964 4544
rect 5052 4536 5060 4544
rect 5548 4536 5556 4544
rect 6124 4536 6132 4544
rect 6188 4536 6196 4544
rect 6348 4536 6356 4544
rect 6364 4536 6372 4544
rect 6396 4536 6404 4544
rect 6428 4536 6436 4544
rect 6444 4536 6452 4544
rect 6492 4536 6500 4544
rect 6748 4536 6756 4544
rect 6828 4536 6836 4544
rect 6940 4536 6948 4544
rect 28 4496 36 4504
rect 92 4496 100 4504
rect 156 4496 164 4504
rect 428 4516 436 4524
rect 492 4516 500 4524
rect 588 4516 596 4524
rect 620 4516 628 4524
rect 668 4516 676 4524
rect 764 4516 772 4524
rect 892 4516 900 4524
rect 940 4516 948 4524
rect 1084 4516 1092 4524
rect 1292 4516 1300 4524
rect 1468 4516 1476 4524
rect 1516 4516 1524 4524
rect 1660 4516 1668 4524
rect 1708 4516 1716 4524
rect 1820 4516 1828 4524
rect 1964 4516 1972 4524
rect 1996 4516 2004 4524
rect 2060 4516 2068 4524
rect 2156 4516 2164 4524
rect 2220 4516 2228 4524
rect 2300 4516 2308 4524
rect 2348 4516 2356 4524
rect 2364 4516 2372 4524
rect 2444 4516 2452 4524
rect 2492 4516 2500 4524
rect 2572 4516 2580 4524
rect 2716 4516 2724 4524
rect 2748 4516 2756 4524
rect 2764 4516 2772 4524
rect 2796 4516 2804 4524
rect 2828 4516 2836 4524
rect 2892 4516 2900 4524
rect 2924 4516 2932 4524
rect 3004 4516 3012 4524
rect 3164 4518 3172 4526
rect 3356 4518 3364 4526
rect 3452 4516 3460 4524
rect 3484 4516 3492 4524
rect 3580 4516 3588 4524
rect 3596 4516 3604 4524
rect 3692 4516 3700 4524
rect 460 4496 468 4504
rect 524 4496 532 4504
rect 572 4496 580 4504
rect 636 4496 644 4504
rect 956 4496 964 4504
rect 1052 4496 1060 4504
rect 1132 4496 1140 4504
rect 1548 4496 1556 4504
rect 1692 4496 1700 4504
rect 1756 4496 1764 4504
rect 1900 4496 1908 4504
rect 1932 4496 1940 4504
rect 2204 4496 2212 4504
rect 2636 4496 2644 4504
rect 3516 4496 3524 4504
rect 3708 4496 3716 4504
rect 3836 4496 3844 4504
rect 3916 4516 3924 4524
rect 3932 4516 3940 4524
rect 4156 4518 4164 4526
rect 4284 4516 4292 4524
rect 4332 4516 4340 4524
rect 4412 4516 4420 4524
rect 4476 4516 4484 4524
rect 4588 4516 4596 4524
rect 4604 4516 4612 4524
rect 4012 4496 4020 4504
rect 4668 4516 4676 4524
rect 4700 4516 4708 4524
rect 4764 4516 4772 4524
rect 4812 4516 4820 4524
rect 4844 4516 4852 4524
rect 4892 4516 4900 4524
rect 4908 4516 4916 4524
rect 4940 4516 4948 4524
rect 4988 4516 4996 4524
rect 5036 4516 5044 4524
rect 5084 4516 5092 4524
rect 5132 4516 5140 4524
rect 5148 4516 5156 4524
rect 5212 4516 5220 4524
rect 5228 4516 5236 4524
rect 5244 4516 5252 4524
rect 5308 4516 5316 4524
rect 5356 4516 5364 4524
rect 5372 4516 5380 4524
rect 5388 4516 5396 4524
rect 5436 4516 5444 4524
rect 5500 4516 5508 4524
rect 5564 4516 5572 4524
rect 5580 4516 5588 4524
rect 5596 4516 5604 4524
rect 5660 4516 5668 4524
rect 5708 4516 5716 4524
rect 5756 4516 5764 4524
rect 5804 4516 5812 4524
rect 5820 4516 5828 4524
rect 5868 4516 5876 4524
rect 5980 4516 5988 4524
rect 6060 4516 6068 4524
rect 6076 4516 6084 4524
rect 6140 4516 6148 4524
rect 6172 4516 6180 4524
rect 6204 4516 6212 4524
rect 6284 4516 6292 4524
rect 6300 4516 6308 4524
rect 6332 4516 6340 4524
rect 6364 4516 6372 4524
rect 6412 4516 6420 4524
rect 4796 4496 4804 4504
rect 5004 4496 5012 4504
rect 5116 4496 5124 4504
rect 6300 4496 6308 4504
rect 6476 4516 6484 4524
rect 6524 4516 6532 4524
rect 6540 4516 6548 4524
rect 6572 4516 6580 4524
rect 6588 4516 6596 4524
rect 6620 4516 6628 4524
rect 6668 4516 6676 4524
rect 6684 4516 6692 4524
rect 6700 4516 6708 4524
rect 6780 4516 6788 4524
rect 6844 4516 6852 4524
rect 6892 4516 6900 4524
rect 6956 4516 6964 4524
rect 7132 4536 7140 4544
rect 7212 4536 7220 4544
rect 7404 4536 7412 4544
rect 7004 4516 7012 4524
rect 7100 4516 7108 4524
rect 7148 4518 7156 4526
rect 6636 4496 6644 4504
rect 364 4476 372 4484
rect 1772 4476 1780 4484
rect 2236 4476 2244 4484
rect 3036 4476 3044 4484
rect 6092 4456 6100 4464
rect 6284 4456 6292 4464
rect 124 4436 132 4444
rect 332 4436 340 4444
rect 556 4436 564 4444
rect 604 4436 612 4444
rect 748 4436 756 4444
rect 876 4436 884 4444
rect 892 4436 900 4444
rect 988 4436 996 4444
rect 1068 4436 1076 4444
rect 1228 4436 1236 4444
rect 1340 4436 1348 4444
rect 2188 4436 2196 4444
rect 2220 4436 2228 4444
rect 2268 4436 2276 4444
rect 2396 4436 2404 4444
rect 2428 4436 2436 4444
rect 2476 4436 2484 4444
rect 2796 4436 2804 4444
rect 3228 4436 3236 4444
rect 3420 4436 3428 4444
rect 4028 4436 4036 4444
rect 5084 4436 5092 4444
rect 5164 4436 5172 4444
rect 5404 4436 5412 4444
rect 5612 4436 5620 4444
rect 5916 4436 5924 4444
rect 1411 4406 1419 4414
rect 1421 4406 1429 4414
rect 1431 4406 1439 4414
rect 1441 4406 1449 4414
rect 1451 4406 1459 4414
rect 1461 4406 1469 4414
rect 4419 4406 4427 4414
rect 4429 4406 4437 4414
rect 4439 4406 4447 4414
rect 4449 4406 4457 4414
rect 4459 4406 4467 4414
rect 4469 4406 4477 4414
rect 156 4376 164 4384
rect 1708 4376 1716 4384
rect 2028 4376 2036 4384
rect 2220 4376 2228 4384
rect 2252 4376 2260 4384
rect 2604 4376 2612 4384
rect 2892 4376 2900 4384
rect 3052 4376 3060 4384
rect 3100 4376 3108 4384
rect 3356 4376 3364 4384
rect 3436 4376 3444 4384
rect 3500 4376 3508 4384
rect 3548 4376 3556 4384
rect 3612 4376 3620 4384
rect 3756 4376 3764 4384
rect 3948 4376 3956 4384
rect 3964 4376 3972 4384
rect 3996 4376 4004 4384
rect 4236 4376 4244 4384
rect 4668 4376 4676 4384
rect 4764 4376 4772 4384
rect 4876 4376 4884 4384
rect 4988 4376 4996 4384
rect 5212 4376 5220 4384
rect 5500 4376 5508 4384
rect 6156 4376 6164 4384
rect 7196 4376 7204 4384
rect 5436 4356 5444 4364
rect 6236 4356 6244 4364
rect 1692 4336 1700 4344
rect 1900 4336 1908 4344
rect 2140 4336 2148 4344
rect 2332 4336 2340 4344
rect 2620 4336 2628 4344
rect 2908 4336 2916 4344
rect 5676 4336 5684 4344
rect 5836 4336 5844 4344
rect 6300 4336 6308 4344
rect 6364 4336 6372 4344
rect 6716 4336 6724 4344
rect 140 4316 148 4324
rect 220 4316 228 4324
rect 620 4316 628 4324
rect 668 4316 676 4324
rect 924 4316 932 4324
rect 364 4296 372 4304
rect 396 4296 404 4304
rect 700 4296 708 4304
rect 748 4296 756 4304
rect 44 4280 52 4288
rect 108 4276 116 4284
rect 172 4276 180 4284
rect 268 4276 276 4284
rect 412 4276 420 4284
rect 492 4276 500 4284
rect 508 4276 516 4284
rect 604 4276 612 4284
rect 652 4276 660 4284
rect 860 4296 868 4304
rect 892 4296 900 4304
rect 924 4296 932 4304
rect 972 4296 980 4304
rect 1052 4316 1060 4324
rect 1148 4316 1156 4324
rect 1324 4316 1332 4324
rect 1564 4316 1572 4324
rect 1084 4296 1092 4304
rect 1180 4296 1188 4304
rect 1228 4296 1236 4304
rect 1372 4296 1380 4304
rect 1420 4296 1428 4304
rect 1532 4296 1540 4304
rect 1724 4316 1732 4324
rect 1612 4296 1620 4304
rect 1708 4296 1716 4304
rect 2076 4316 2084 4324
rect 2172 4316 2180 4324
rect 2284 4316 2292 4324
rect 2300 4316 2308 4324
rect 2380 4316 2388 4324
rect 2396 4316 2404 4324
rect 2508 4316 2516 4324
rect 2524 4316 2532 4324
rect 2588 4316 2596 4324
rect 2732 4316 2740 4324
rect 2876 4316 2884 4324
rect 3292 4316 3300 4324
rect 3452 4316 3460 4324
rect 3532 4316 3540 4324
rect 3644 4316 3652 4324
rect 5772 4316 5780 4324
rect 1788 4296 1796 4304
rect 1980 4296 1988 4304
rect 2060 4296 2068 4304
rect 2156 4296 2164 4304
rect 2188 4296 2196 4304
rect 2252 4296 2260 4304
rect 2316 4296 2324 4304
rect 2412 4296 2420 4304
rect 2572 4296 2580 4304
rect 2604 4296 2612 4304
rect 2652 4296 2660 4304
rect 2700 4296 2708 4304
rect 2796 4296 2804 4304
rect 2892 4296 2900 4304
rect 3004 4296 3012 4304
rect 3084 4296 3092 4304
rect 3228 4294 3236 4302
rect 3308 4296 3316 4304
rect 3324 4296 3332 4304
rect 3388 4296 3396 4304
rect 3404 4296 3412 4304
rect 3500 4296 3508 4304
rect 3580 4296 3588 4304
rect 3612 4296 3620 4304
rect 3692 4296 3700 4304
rect 3724 4296 3732 4304
rect 3836 4296 3844 4304
rect 3884 4296 3892 4304
rect 4156 4294 4164 4302
rect 4508 4296 4516 4304
rect 4620 4296 4628 4304
rect 4636 4296 4644 4304
rect 4732 4296 4740 4304
rect 4780 4296 4788 4304
rect 4796 4296 4804 4304
rect 4812 4296 4820 4304
rect 4892 4296 4900 4304
rect 5004 4296 5012 4304
rect 5020 4296 5028 4304
rect 5068 4296 5076 4304
rect 5084 4296 5092 4304
rect 5116 4296 5124 4304
rect 5148 4296 5156 4304
rect 5196 4296 5204 4304
rect 5244 4296 5252 4304
rect 5260 4296 5268 4304
rect 5292 4296 5300 4304
rect 5324 4296 5332 4304
rect 5356 4296 5364 4304
rect 5420 4296 5428 4304
rect 5468 4296 5476 4304
rect 5484 4296 5492 4304
rect 5532 4296 5540 4304
rect 5564 4296 5572 4304
rect 5596 4296 5604 4304
rect 5612 4296 5620 4304
rect 860 4276 868 4284
rect 876 4276 884 4284
rect 908 4276 916 4284
rect 988 4276 996 4284
rect 1004 4276 1012 4284
rect 1180 4276 1188 4284
rect 1292 4276 1300 4284
rect 1372 4276 1380 4284
rect 1436 4276 1444 4284
rect 1500 4276 1508 4284
rect 1628 4276 1636 4284
rect 1740 4276 1748 4284
rect 1868 4276 1876 4284
rect 1932 4276 1940 4284
rect 2236 4276 2244 4284
rect 2364 4276 2372 4284
rect 2428 4276 2436 4284
rect 2476 4276 2484 4284
rect 2508 4276 2516 4284
rect 2572 4276 2580 4284
rect 2684 4276 2692 4284
rect 2780 4276 2788 4284
rect 3212 4276 3220 4284
rect 3484 4276 3492 4284
rect 3596 4276 3604 4284
rect 3708 4276 3716 4284
rect 4348 4276 4356 4284
rect 4444 4276 4452 4284
rect 4492 4276 4500 4284
rect 4844 4276 4852 4284
rect 4892 4276 4900 4284
rect 4956 4276 4964 4284
rect 4988 4276 4996 4284
rect 5100 4276 5108 4284
rect 5132 4276 5140 4284
rect 5180 4276 5188 4284
rect 5276 4276 5284 4284
rect 5340 4276 5348 4284
rect 5548 4276 5556 4284
rect 5612 4276 5620 4284
rect 124 4256 132 4264
rect 140 4256 148 4264
rect 220 4256 228 4264
rect 236 4256 244 4264
rect 316 4256 324 4264
rect 348 4256 356 4264
rect 428 4256 436 4264
rect 748 4256 756 4264
rect 1132 4256 1140 4264
rect 1308 4256 1316 4264
rect 1660 4256 1668 4264
rect 1820 4256 1828 4264
rect 1916 4256 1924 4264
rect 2012 4256 2020 4264
rect 2348 4256 2356 4264
rect 2460 4256 2468 4264
rect 2668 4256 2676 4264
rect 2748 4256 2756 4264
rect 3468 4256 3476 4264
rect 3980 4256 3988 4264
rect 4012 4256 4020 4264
rect 4156 4256 4164 4264
rect 4940 4256 4948 4264
rect 5324 4256 5332 4264
rect 5388 4256 5396 4264
rect 5564 4256 5572 4264
rect 5708 4296 5716 4304
rect 5740 4296 5748 4304
rect 5756 4296 5764 4304
rect 5804 4296 5812 4304
rect 5884 4296 5892 4304
rect 6044 4296 6052 4304
rect 6172 4296 6180 4304
rect 6268 4296 6276 4304
rect 6588 4316 6596 4324
rect 6332 4296 6340 4304
rect 6748 4316 6756 4324
rect 6492 4294 6500 4302
rect 6636 4296 6644 4304
rect 6668 4296 6676 4304
rect 6780 4296 6788 4304
rect 6796 4296 6804 4304
rect 6892 4316 6900 4324
rect 7180 4316 7188 4324
rect 7052 4296 7060 4304
rect 7148 4296 7156 4304
rect 7180 4296 7188 4304
rect 7308 4296 7316 4304
rect 5724 4276 5732 4284
rect 5788 4276 5796 4284
rect 5868 4276 5876 4284
rect 5900 4276 5908 4284
rect 6220 4276 6228 4284
rect 6284 4276 6292 4284
rect 6348 4276 6356 4284
rect 6524 4276 6532 4284
rect 6556 4276 6564 4284
rect 6588 4276 6596 4284
rect 6652 4276 6660 4284
rect 6716 4276 6724 4284
rect 6812 4276 6820 4284
rect 6828 4276 6836 4284
rect 6924 4276 6932 4284
rect 7052 4276 7060 4284
rect 7100 4276 7108 4284
rect 7132 4276 7140 4284
rect 7292 4276 7300 4284
rect 5644 4256 5652 4264
rect 6028 4256 6036 4264
rect 6204 4256 6212 4264
rect 6300 4256 6308 4264
rect 12 4236 20 4244
rect 252 4236 260 4244
rect 460 4236 468 4244
rect 540 4236 548 4244
rect 620 4236 628 4244
rect 668 4236 676 4244
rect 828 4236 836 4244
rect 1036 4236 1044 4244
rect 1196 4236 1204 4244
rect 1324 4236 1332 4244
rect 1388 4236 1396 4244
rect 1580 4236 1588 4244
rect 1644 4236 1652 4244
rect 1756 4236 1764 4244
rect 1804 4236 1812 4244
rect 1836 4236 1844 4244
rect 2092 4236 2100 4244
rect 2220 4236 2228 4244
rect 2444 4236 2452 4244
rect 2492 4236 2500 4244
rect 2732 4236 2740 4244
rect 2780 4236 2788 4244
rect 3036 4236 3044 4244
rect 3052 4236 3060 4244
rect 3100 4236 3108 4244
rect 3660 4236 3668 4244
rect 3756 4236 3764 4244
rect 4028 4236 4036 4244
rect 4604 4236 4612 4244
rect 5372 4236 5380 4244
rect 6876 4236 6884 4244
rect 6940 4236 6948 4244
rect 2915 4206 2923 4214
rect 2925 4206 2933 4214
rect 2935 4206 2943 4214
rect 2945 4206 2953 4214
rect 2955 4206 2963 4214
rect 2965 4206 2973 4214
rect 5923 4206 5931 4214
rect 5933 4206 5941 4214
rect 5943 4206 5951 4214
rect 5953 4206 5961 4214
rect 5963 4206 5971 4214
rect 5973 4206 5981 4214
rect 460 4176 468 4184
rect 700 4176 708 4184
rect 1628 4176 1636 4184
rect 2156 4176 2164 4184
rect 2268 4176 2276 4184
rect 2300 4176 2308 4184
rect 2460 4176 2468 4184
rect 2636 4176 2644 4184
rect 2716 4176 2724 4184
rect 2892 4176 2900 4184
rect 3020 4176 3028 4184
rect 3260 4176 3268 4184
rect 3340 4176 3348 4184
rect 3788 4176 3796 4184
rect 3836 4176 3844 4184
rect 4076 4176 4084 4184
rect 4172 4176 4180 4184
rect 4236 4176 4244 4184
rect 4508 4176 4516 4184
rect 4588 4176 4596 4184
rect 4828 4176 4836 4184
rect 5180 4176 5188 4184
rect 5196 4176 5204 4184
rect 5356 4176 5364 4184
rect 6908 4176 6916 4184
rect 6972 4176 6980 4184
rect 156 4156 164 4164
rect 364 4156 372 4164
rect 380 4156 388 4164
rect 620 4156 628 4164
rect 860 4156 868 4164
rect 940 4156 948 4164
rect 1020 4156 1028 4164
rect 1116 4156 1124 4164
rect 1260 4156 1268 4164
rect 1372 4156 1380 4164
rect 1404 4156 1412 4164
rect 1500 4156 1508 4164
rect 1820 4156 1828 4164
rect 1980 4156 1988 4164
rect 2108 4156 2116 4164
rect 2188 4156 2196 4164
rect 2236 4156 2244 4164
rect 2252 4156 2260 4164
rect 2620 4156 2628 4164
rect 2828 4156 2836 4164
rect 2844 4156 2852 4164
rect 3676 4156 3684 4164
rect 4572 4156 4580 4164
rect 4924 4156 4932 4164
rect 108 4136 116 4144
rect 428 4136 436 4144
rect 524 4136 532 4144
rect 604 4136 612 4144
rect 636 4136 644 4144
rect 732 4136 740 4144
rect 812 4136 820 4144
rect 1276 4136 1284 4144
rect 1308 4136 1316 4144
rect 1532 4136 1540 4144
rect 1580 4136 1588 4144
rect 1596 4136 1604 4144
rect 1708 4136 1716 4144
rect 1772 4136 1780 4144
rect 1900 4136 1908 4144
rect 2316 4136 2324 4144
rect 2348 4136 2356 4144
rect 2380 4136 2388 4144
rect 2428 4136 2436 4144
rect 2460 4136 2468 4144
rect 2476 4136 2484 4144
rect 2524 4136 2532 4144
rect 2556 4136 2564 4144
rect 2572 4136 2580 4144
rect 2652 4136 2660 4144
rect 44 4116 52 4124
rect 76 4116 84 4124
rect 204 4116 212 4124
rect 220 4116 228 4124
rect 284 4116 292 4124
rect 412 4116 420 4124
rect 780 4116 788 4124
rect 796 4116 804 4124
rect 844 4116 852 4124
rect 892 4116 900 4124
rect 956 4116 964 4124
rect 972 4116 980 4124
rect 1020 4116 1028 4124
rect 1036 4116 1044 4124
rect 1068 4116 1076 4124
rect 1180 4116 1188 4124
rect 1228 4116 1236 4124
rect 1340 4116 1348 4124
rect 1372 4116 1380 4124
rect 1580 4116 1588 4124
rect 1692 4116 1700 4124
rect 60 4096 68 4104
rect 140 4096 148 4104
rect 236 4096 244 4104
rect 252 4096 260 4104
rect 1004 4096 1012 4104
rect 1052 4096 1060 4104
rect 1324 4096 1332 4104
rect 1740 4096 1748 4104
rect 1804 4116 1812 4124
rect 1852 4116 1860 4124
rect 1932 4116 1940 4124
rect 1948 4116 1956 4124
rect 1996 4116 2004 4124
rect 2076 4116 2084 4124
rect 2124 4116 2132 4124
rect 2732 4136 2740 4144
rect 2764 4136 2772 4144
rect 2796 4136 2804 4144
rect 2828 4136 2836 4144
rect 2908 4136 2916 4144
rect 3084 4136 3092 4144
rect 3180 4136 3188 4144
rect 2396 4116 2404 4124
rect 2412 4116 2420 4124
rect 2476 4116 2484 4124
rect 2508 4116 2516 4124
rect 2540 4116 2548 4124
rect 2668 4116 2676 4124
rect 2236 4096 2244 4104
rect 2284 4096 2292 4104
rect 2604 4096 2612 4104
rect 2748 4116 2756 4124
rect 2780 4116 2788 4124
rect 2812 4116 2820 4124
rect 2988 4116 2996 4124
rect 3068 4116 3076 4124
rect 3292 4136 3300 4144
rect 3388 4136 3396 4144
rect 3452 4136 3460 4144
rect 3516 4136 3524 4144
rect 3548 4136 3556 4144
rect 3676 4136 3684 4144
rect 3708 4136 3716 4144
rect 3724 4136 3732 4144
rect 3884 4136 3892 4144
rect 3964 4136 3972 4144
rect 4060 4136 4068 4144
rect 4092 4136 4100 4144
rect 4188 4136 4196 4144
rect 4348 4136 4356 4144
rect 4396 4136 4404 4144
rect 4492 4136 4500 4144
rect 4748 4136 4756 4144
rect 4780 4136 4788 4144
rect 4876 4136 4884 4144
rect 5772 4156 5780 4164
rect 6028 4156 6036 4164
rect 6156 4156 6164 4164
rect 6300 4156 6308 4164
rect 6812 4156 6820 4164
rect 7292 4156 7300 4164
rect 4972 4136 4980 4144
rect 5020 4136 5028 4144
rect 5260 4136 5268 4144
rect 5292 4136 5300 4144
rect 5564 4136 5572 4144
rect 5596 4136 5604 4144
rect 5708 4136 5716 4144
rect 5772 4136 5780 4144
rect 5820 4136 5828 4144
rect 5852 4136 5860 4144
rect 5884 4136 5892 4144
rect 5900 4136 5908 4144
rect 6012 4136 6020 4144
rect 6076 4136 6084 4144
rect 6140 4136 6148 4144
rect 6204 4136 6212 4144
rect 6316 4136 6324 4144
rect 6348 4136 6356 4144
rect 6380 4136 6388 4144
rect 6412 4136 6420 4144
rect 6444 4136 6452 4144
rect 6460 4136 6468 4144
rect 6572 4136 6580 4144
rect 6652 4136 6660 4144
rect 6748 4136 6756 4144
rect 3228 4096 3236 4104
rect 3244 4096 3252 4104
rect 3324 4096 3332 4104
rect 3372 4116 3380 4124
rect 3436 4116 3444 4124
rect 3468 4116 3476 4124
rect 3564 4116 3572 4124
rect 3612 4116 3620 4124
rect 3628 4116 3636 4124
rect 3724 4116 3732 4124
rect 3820 4116 3828 4124
rect 3868 4116 3876 4124
rect 3996 4116 4004 4124
rect 4108 4116 4116 4124
rect 4204 4116 4212 4124
rect 4476 4116 4484 4124
rect 4540 4116 4548 4124
rect 4652 4116 4660 4124
rect 4716 4118 4724 4126
rect 3500 4096 3508 4104
rect 3740 4096 3748 4104
rect 4140 4096 4148 4104
rect 4812 4096 4820 4104
rect 4860 4116 4868 4124
rect 4892 4116 4900 4124
rect 4956 4116 4964 4124
rect 4988 4116 4996 4124
rect 5052 4118 5060 4126
rect 5228 4116 5236 4124
rect 5276 4116 5284 4124
rect 5340 4116 5348 4124
rect 5388 4116 5396 4124
rect 5516 4116 5524 4124
rect 5612 4116 5620 4124
rect 5244 4096 5252 4104
rect 5692 4116 5700 4124
rect 5724 4116 5732 4124
rect 5772 4116 5780 4124
rect 5804 4116 5812 4124
rect 5836 4116 5844 4124
rect 5868 4116 5876 4124
rect 5660 4096 5668 4104
rect 5932 4116 5940 4124
rect 6044 4116 6052 4124
rect 6060 4116 6068 4124
rect 6092 4116 6100 4124
rect 6124 4116 6132 4124
rect 6188 4116 6196 4124
rect 6220 4116 6228 4124
rect 6268 4116 6276 4124
rect 6364 4116 6372 4124
rect 6428 4116 6436 4124
rect 6476 4116 6484 4124
rect 6396 4096 6404 4104
rect 6556 4116 6564 4124
rect 6700 4116 6708 4124
rect 6780 4116 6788 4124
rect 6796 4116 6804 4124
rect 6892 4116 6900 4124
rect 6940 4116 6948 4124
rect 6956 4116 6964 4124
rect 7052 4116 7060 4124
rect 7084 4116 7092 4124
rect 7228 4116 7236 4124
rect 7260 4116 7268 4124
rect 6556 4096 6564 4104
rect 28 4076 36 4084
rect 556 4076 564 4084
rect 1084 4076 1092 4084
rect 1116 4076 1124 4084
rect 2572 4076 2580 4084
rect 3036 4076 3044 4084
rect 5308 4076 5316 4084
rect 5404 4076 5412 4084
rect 6508 4076 6516 4084
rect 6588 4076 6596 4084
rect 7164 4076 7172 4084
rect 2028 4056 2036 4064
rect 5612 4056 5620 4064
rect 6092 4056 6100 4064
rect 6252 4056 6260 4064
rect 44 4036 52 4044
rect 124 4036 132 4044
rect 284 4036 292 4044
rect 396 4036 404 4044
rect 748 4036 756 4044
rect 1068 4036 1076 4044
rect 1148 4036 1156 4044
rect 1196 4036 1204 4044
rect 1372 4036 1380 4044
rect 1564 4036 1572 4044
rect 2044 4036 2052 4044
rect 2380 4036 2388 4044
rect 3212 4036 3220 4044
rect 3676 4036 3684 4044
rect 5196 4036 5204 4044
rect 1411 4006 1419 4014
rect 1421 4006 1429 4014
rect 1431 4006 1439 4014
rect 1441 4006 1449 4014
rect 1451 4006 1459 4014
rect 1461 4006 1469 4014
rect 4419 4006 4427 4014
rect 4429 4006 4437 4014
rect 4439 4006 4447 4014
rect 4449 4006 4457 4014
rect 4459 4006 4467 4014
rect 4469 4006 4477 4014
rect 92 3976 100 3984
rect 236 3976 244 3984
rect 1100 3976 1108 3984
rect 2028 3976 2036 3984
rect 3468 3976 3476 3984
rect 3948 3976 3956 3984
rect 3996 3976 4004 3984
rect 4284 3976 4292 3984
rect 4908 3976 4916 3984
rect 5532 3976 5540 3984
rect 6060 3976 6068 3984
rect 6252 3976 6260 3984
rect 6300 3976 6308 3984
rect 6156 3956 6164 3964
rect 6684 3956 6692 3964
rect 1948 3936 1956 3944
rect 4316 3936 4324 3944
rect 5052 3936 5060 3944
rect 5116 3936 5124 3944
rect 5260 3936 5268 3944
rect 5292 3936 5300 3944
rect 6380 3936 6388 3944
rect 6508 3936 6516 3944
rect 6860 3936 6868 3944
rect 7148 3936 7156 3944
rect 7196 3936 7204 3944
rect 7228 3936 7236 3944
rect 44 3916 52 3924
rect 60 3916 68 3924
rect 348 3916 356 3924
rect 476 3916 484 3924
rect 540 3916 548 3924
rect 572 3916 580 3924
rect 652 3916 660 3924
rect 700 3916 708 3924
rect 780 3916 788 3924
rect 812 3916 820 3924
rect 1036 3916 1044 3924
rect 1084 3916 1092 3924
rect 92 3896 100 3904
rect 284 3896 292 3904
rect 316 3896 324 3904
rect 460 3896 468 3904
rect 876 3896 884 3904
rect 1180 3896 1188 3904
rect 1196 3896 1204 3904
rect 1212 3896 1220 3904
rect 1276 3896 1284 3904
rect 1692 3896 1700 3904
rect 1820 3896 1828 3904
rect 1884 3896 1892 3904
rect 1932 3896 1940 3904
rect 1980 3896 1988 3904
rect 1996 3896 2004 3904
rect 2060 3896 2068 3904
rect 2188 3896 2196 3904
rect 2236 3896 2244 3904
rect 2284 3896 2292 3904
rect 2364 3896 2372 3904
rect 2444 3916 2452 3924
rect 2716 3916 2724 3924
rect 2876 3916 2884 3924
rect 3036 3916 3044 3924
rect 3820 3916 3828 3924
rect 3916 3916 3924 3924
rect 3980 3916 3988 3924
rect 4108 3916 4116 3924
rect 4172 3916 4180 3924
rect 4188 3916 4196 3924
rect 4268 3916 4276 3924
rect 5228 3916 5236 3924
rect 5516 3916 5524 3924
rect 5756 3916 5764 3924
rect 2476 3896 2484 3904
rect 2620 3896 2628 3904
rect 2700 3896 2708 3904
rect 3084 3896 3092 3904
rect 3132 3896 3140 3904
rect 3196 3896 3204 3904
rect 3308 3896 3316 3904
rect 3596 3894 3604 3902
rect 3724 3896 3732 3904
rect 3884 3896 3892 3904
rect 4076 3896 4084 3904
rect 4140 3896 4148 3904
rect 4412 3894 4420 3902
rect 4668 3894 4676 3902
rect 4732 3896 4740 3904
rect 4796 3896 4804 3904
rect 4844 3896 4852 3904
rect 4860 3896 4868 3904
rect 4892 3896 4900 3904
rect 4940 3896 4948 3904
rect 4956 3896 4964 3904
rect 4988 3896 4996 3904
rect 5036 3896 5044 3904
rect 5052 3896 5060 3904
rect 5116 3896 5124 3904
rect 5212 3896 5220 3904
rect 5260 3896 5268 3904
rect 5884 3916 5892 3924
rect 6108 3916 6116 3924
rect 6444 3916 6452 3924
rect 6780 3916 6788 3924
rect 5420 3894 5428 3902
rect 5660 3894 5668 3902
rect 5804 3896 5812 3904
rect 5852 3896 5860 3904
rect 12 3876 20 3884
rect 108 3876 116 3884
rect 124 3876 132 3884
rect 268 3876 276 3884
rect 300 3876 308 3884
rect 364 3876 372 3884
rect 460 3876 468 3884
rect 524 3876 532 3884
rect 572 3876 580 3884
rect 620 3876 628 3884
rect 684 3876 692 3884
rect 716 3876 724 3884
rect 764 3876 772 3884
rect 812 3876 820 3884
rect 860 3876 868 3884
rect 924 3876 932 3884
rect 1020 3876 1028 3884
rect 1068 3876 1076 3884
rect 1116 3876 1124 3884
rect 1260 3876 1268 3884
rect 1388 3876 1396 3884
rect 1404 3876 1412 3884
rect 1564 3876 1572 3884
rect 1580 3876 1588 3884
rect 1676 3876 1684 3884
rect 236 3856 244 3864
rect 540 3856 548 3864
rect 636 3856 644 3864
rect 652 3856 660 3864
rect 716 3856 724 3864
rect 732 3856 740 3864
rect 844 3856 852 3864
rect 1132 3856 1140 3864
rect 1212 3856 1220 3864
rect 1724 3856 1732 3864
rect 1836 3876 1844 3884
rect 1900 3876 1908 3884
rect 2204 3876 2212 3884
rect 2380 3876 2388 3884
rect 2396 3876 2404 3884
rect 2492 3876 2500 3884
rect 2508 3876 2516 3884
rect 2604 3876 2612 3884
rect 2652 3876 2660 3884
rect 2716 3876 2724 3884
rect 2764 3876 2772 3884
rect 2844 3876 2852 3884
rect 2924 3876 2932 3884
rect 3004 3876 3012 3884
rect 3052 3876 3060 3884
rect 3148 3876 3156 3884
rect 3212 3876 3220 3884
rect 3324 3876 3332 3884
rect 2140 3856 2148 3864
rect 2284 3856 2292 3864
rect 2316 3856 2324 3864
rect 2860 3856 2868 3864
rect 2988 3856 2996 3864
rect 3164 3856 3172 3864
rect 3260 3856 3268 3864
rect 3324 3856 3332 3864
rect 3436 3876 3444 3884
rect 3564 3876 3572 3884
rect 3852 3876 3860 3884
rect 3868 3876 3876 3884
rect 3932 3876 3940 3884
rect 4028 3880 4036 3888
rect 4044 3876 4052 3884
rect 4060 3876 4068 3884
rect 4156 3876 4164 3884
rect 4236 3876 4244 3884
rect 4780 3876 4788 3884
rect 4972 3876 4980 3884
rect 5036 3876 5044 3884
rect 5100 3876 5108 3884
rect 5164 3876 5172 3884
rect 5276 3876 5284 3884
rect 5452 3876 5460 3884
rect 5484 3876 5492 3884
rect 5692 3876 5700 3884
rect 5724 3876 5732 3884
rect 5772 3876 5780 3884
rect 5820 3876 5828 3884
rect 5836 3876 5844 3884
rect 5900 3876 5908 3884
rect 5980 3896 5988 3904
rect 6028 3896 6036 3904
rect 6140 3896 6148 3904
rect 6188 3896 6196 3904
rect 6204 3896 6212 3904
rect 6220 3896 6228 3904
rect 6284 3896 6292 3904
rect 6332 3896 6340 3904
rect 6348 3896 6356 3904
rect 6380 3896 6388 3904
rect 6412 3896 6420 3904
rect 6492 3896 6500 3904
rect 6508 3896 6516 3904
rect 6572 3896 6580 3904
rect 6620 3896 6628 3904
rect 6636 3896 6644 3904
rect 6652 3896 6660 3904
rect 6668 3896 6676 3904
rect 6828 3916 6836 3924
rect 7180 3916 7188 3924
rect 6076 3876 6084 3884
rect 6364 3876 6372 3884
rect 6492 3876 6500 3884
rect 6572 3876 6580 3884
rect 6828 3896 6836 3904
rect 6972 3896 6980 3904
rect 7084 3896 7092 3904
rect 7100 3896 7108 3904
rect 7260 3896 7268 3904
rect 7276 3896 7284 3904
rect 6748 3876 6756 3884
rect 6844 3876 6852 3884
rect 7020 3876 7028 3884
rect 7052 3876 7060 3884
rect 7148 3876 7156 3884
rect 3452 3856 3460 3864
rect 3756 3856 3764 3864
rect 3804 3856 3812 3864
rect 4316 3856 4324 3864
rect 4412 3856 4420 3864
rect 4668 3856 4676 3864
rect 4764 3856 4772 3864
rect 5084 3856 5092 3864
rect 5180 3856 5188 3864
rect 6012 3856 6020 3864
rect 6540 3856 6548 3864
rect 7052 3856 7060 3864
rect 44 3836 52 3844
rect 188 3836 196 3844
rect 348 3836 356 3844
rect 412 3836 420 3844
rect 908 3836 916 3844
rect 988 3836 996 3844
rect 1036 3836 1044 3844
rect 1244 3836 1252 3844
rect 1324 3836 1332 3844
rect 1532 3836 1540 3844
rect 1612 3836 1620 3844
rect 1756 3836 1764 3844
rect 2124 3836 2132 3844
rect 2156 3836 2164 3844
rect 2268 3836 2276 3844
rect 2332 3836 2340 3844
rect 2428 3836 2436 3844
rect 2572 3836 2580 3844
rect 2668 3836 2676 3844
rect 2732 3836 2740 3844
rect 2780 3836 2788 3844
rect 2876 3836 2884 3844
rect 3100 3836 3108 3844
rect 3324 3836 3332 3844
rect 3420 3836 3428 3844
rect 3740 3836 3748 3844
rect 3836 3836 3844 3844
rect 4204 3836 4212 3844
rect 4268 3836 4276 3844
rect 4540 3836 4548 3844
rect 4748 3836 4756 3844
rect 4988 3836 4996 3844
rect 5500 3836 5508 3844
rect 6092 3836 6100 3844
rect 7068 3836 7076 3844
rect 7180 3836 7188 3844
rect 2915 3806 2923 3814
rect 2925 3806 2933 3814
rect 2935 3806 2943 3814
rect 2945 3806 2953 3814
rect 2955 3806 2963 3814
rect 2965 3806 2973 3814
rect 5923 3806 5931 3814
rect 5933 3806 5941 3814
rect 5943 3806 5951 3814
rect 5953 3806 5961 3814
rect 5963 3806 5971 3814
rect 5973 3806 5981 3814
rect 508 3796 516 3804
rect 620 3796 628 3804
rect 956 3796 964 3804
rect 1772 3796 1780 3804
rect 2172 3796 2180 3804
rect 2412 3796 2420 3804
rect 92 3776 100 3784
rect 188 3776 196 3784
rect 252 3776 260 3784
rect 1724 3776 1732 3784
rect 3100 3776 3108 3784
rect 3500 3776 3508 3784
rect 3660 3776 3668 3784
rect 3788 3776 3796 3784
rect 3996 3776 4004 3784
rect 4140 3776 4148 3784
rect 4252 3776 4260 3784
rect 4428 3776 4436 3784
rect 4588 3776 4596 3784
rect 4684 3776 4692 3784
rect 4892 3776 4900 3784
rect 5276 3776 5284 3784
rect 5420 3776 5428 3784
rect 5484 3776 5492 3784
rect 5532 3776 5540 3784
rect 5596 3776 5604 3784
rect 5756 3776 5764 3784
rect 5948 3776 5956 3784
rect 6108 3776 6116 3784
rect 6412 3776 6420 3784
rect 6460 3776 6468 3784
rect 6492 3776 6500 3784
rect 6908 3776 6916 3784
rect 7228 3776 7236 3784
rect 7292 3776 7300 3784
rect 12 3756 20 3764
rect 60 3756 68 3764
rect 220 3756 228 3764
rect 268 3756 276 3764
rect 460 3756 468 3764
rect 476 3756 484 3764
rect 508 3756 516 3764
rect 620 3756 628 3764
rect 780 3756 788 3764
rect 956 3756 964 3764
rect 1324 3756 1332 3764
rect 1772 3756 1780 3764
rect 1948 3756 1956 3764
rect 108 3736 116 3744
rect 140 3736 148 3744
rect 284 3736 292 3744
rect 396 3736 404 3744
rect 428 3736 436 3744
rect 604 3736 612 3744
rect 716 3736 724 3744
rect 764 3736 772 3744
rect 844 3736 852 3744
rect 860 3736 868 3744
rect 892 3736 900 3744
rect 972 3736 980 3744
rect 1068 3736 1076 3744
rect 1084 3736 1092 3744
rect 1180 3736 1188 3744
rect 1676 3736 1684 3744
rect 1980 3756 1988 3764
rect 1996 3756 2004 3764
rect 2108 3756 2116 3764
rect 2172 3756 2180 3764
rect 2204 3756 2212 3764
rect 2268 3756 2276 3764
rect 2412 3756 2420 3764
rect 2444 3756 2452 3764
rect 2860 3756 2868 3764
rect 2876 3756 2884 3764
rect 3004 3756 3012 3764
rect 3356 3756 3364 3764
rect 3676 3756 3684 3764
rect 3804 3756 3812 3764
rect 3836 3756 3844 3764
rect 3852 3756 3860 3764
rect 4172 3756 4180 3764
rect 4220 3756 4228 3764
rect 4444 3756 4452 3764
rect 4524 3756 4532 3764
rect 4700 3756 4708 3764
rect 5116 3756 5124 3764
rect 5292 3756 5300 3764
rect 6556 3756 6564 3764
rect 6700 3756 6708 3764
rect 7340 3756 7348 3764
rect 2012 3736 2020 3744
rect 2252 3736 2260 3744
rect 2316 3736 2324 3744
rect 2412 3736 2420 3744
rect 2460 3736 2468 3744
rect 2556 3736 2564 3744
rect 2604 3736 2612 3744
rect 2620 3736 2628 3744
rect 2716 3736 2724 3744
rect 2748 3736 2756 3744
rect 2780 3736 2788 3744
rect 2812 3736 2820 3744
rect 2844 3736 2852 3744
rect 2908 3736 2916 3744
rect 3260 3736 3268 3744
rect 3292 3736 3300 3744
rect 3356 3736 3364 3744
rect 3388 3736 3396 3744
rect 3500 3736 3508 3744
rect 3532 3736 3540 3744
rect 3644 3736 3652 3744
rect 3708 3736 3716 3744
rect 3740 3736 3748 3744
rect 3900 3736 3908 3744
rect 3996 3736 4004 3744
rect 4028 3736 4036 3744
rect 4156 3736 4164 3744
rect 4252 3736 4260 3744
rect 4300 3736 4308 3744
rect 4332 3736 4340 3744
rect 4348 3736 4356 3744
rect 4364 3736 4372 3744
rect 4412 3736 4420 3744
rect 4572 3736 4580 3744
rect 4636 3736 4644 3744
rect 4652 3736 4660 3744
rect 4732 3736 4740 3744
rect 4908 3736 4916 3744
rect 4940 3736 4948 3744
rect 5020 3736 5028 3744
rect 5036 3736 5044 3744
rect 5068 3736 5076 3744
rect 5100 3736 5108 3744
rect 5212 3736 5220 3744
rect 5340 3736 5348 3744
rect 5404 3736 5412 3744
rect 5468 3736 5476 3744
rect 5580 3736 5588 3744
rect 5644 3736 5652 3744
rect 5676 3736 5684 3744
rect 5692 3736 5700 3744
rect 5740 3736 5748 3744
rect 5884 3736 5892 3744
rect 6060 3736 6068 3744
rect 6172 3736 6180 3744
rect 6284 3736 6292 3744
rect 6476 3736 6484 3744
rect 6540 3736 6548 3744
rect 6604 3736 6612 3744
rect 6716 3736 6724 3744
rect 6844 3736 6852 3744
rect 7052 3736 7060 3744
rect 7116 3736 7124 3744
rect 7180 3736 7188 3744
rect 156 3716 164 3724
rect 236 3716 244 3724
rect 508 3716 516 3724
rect 556 3716 564 3724
rect 588 3716 596 3724
rect 668 3716 676 3724
rect 716 3716 724 3724
rect 828 3716 836 3724
rect 876 3716 884 3724
rect 908 3716 916 3724
rect 1228 3716 1236 3724
rect 1276 3716 1284 3724
rect 1372 3716 1380 3724
rect 1516 3716 1524 3724
rect 1580 3716 1588 3724
rect 1644 3716 1652 3724
rect 1692 3716 1700 3724
rect 1724 3716 1732 3724
rect 1820 3716 1828 3724
rect 1884 3716 1892 3724
rect 1916 3716 1924 3724
rect 1996 3716 2004 3724
rect 2140 3716 2148 3724
rect 2204 3716 2212 3724
rect 2236 3716 2244 3724
rect 2300 3716 2308 3724
rect 2332 3716 2340 3724
rect 2348 3716 2356 3724
rect 2364 3716 2372 3724
rect 2732 3716 2740 3724
rect 2796 3716 2804 3724
rect 3036 3716 3044 3724
rect 3084 3716 3092 3724
rect 3228 3718 3236 3726
rect 3308 3716 3316 3724
rect 3340 3716 3348 3724
rect 3404 3716 3412 3724
rect 3452 3716 3460 3724
rect 3548 3716 3556 3724
rect 3596 3716 3604 3724
rect 3628 3716 3636 3724
rect 3692 3716 3700 3724
rect 3756 3716 3764 3724
rect 3772 3716 3780 3724
rect 3804 3716 3812 3724
rect 3884 3716 3892 3724
rect 3932 3716 3940 3724
rect 3980 3716 3988 3724
rect 4044 3716 4052 3724
rect 4092 3716 4100 3724
rect 4124 3716 4132 3724
rect 4236 3716 4244 3724
rect 4300 3716 4308 3724
rect 4316 3716 4324 3724
rect 4380 3716 4388 3724
rect 4396 3716 4404 3724
rect 4556 3716 4564 3724
rect 4620 3716 4628 3724
rect 4652 3716 4660 3724
rect 4780 3716 4788 3724
rect 4924 3716 4932 3724
rect 396 3696 404 3704
rect 428 3696 436 3704
rect 1244 3696 1252 3704
rect 1260 3696 1268 3704
rect 1356 3696 1364 3704
rect 1532 3696 1540 3704
rect 1596 3696 1604 3704
rect 1660 3696 1668 3704
rect 1836 3696 1844 3704
rect 1900 3696 1908 3704
rect 2572 3696 2580 3704
rect 3340 3696 3348 3704
rect 3468 3696 3476 3704
rect 3596 3696 3604 3704
rect 3708 3696 3716 3704
rect 3852 3696 3860 3704
rect 3916 3696 3924 3704
rect 4108 3696 4116 3704
rect 4476 3696 4484 3704
rect 4588 3696 4596 3704
rect 5004 3716 5012 3724
rect 5052 3716 5060 3724
rect 5148 3716 5156 3724
rect 5180 3716 5188 3724
rect 5228 3716 5236 3724
rect 5244 3716 5252 3724
rect 5324 3716 5332 3724
rect 5340 3716 5348 3724
rect 5388 3716 5396 3724
rect 5452 3716 5460 3724
rect 5516 3716 5524 3724
rect 5564 3716 5572 3724
rect 5644 3716 5652 3724
rect 4972 3696 4980 3704
rect 5164 3696 5172 3704
rect 5276 3696 5284 3704
rect 5420 3696 5428 3704
rect 5532 3696 5540 3704
rect 5708 3716 5716 3724
rect 5868 3716 5876 3724
rect 6060 3716 6068 3724
rect 6076 3716 6084 3724
rect 6156 3716 6164 3724
rect 6188 3716 6196 3724
rect 6300 3716 6308 3724
rect 6428 3716 6436 3724
rect 6492 3716 6500 3724
rect 6588 3716 6596 3724
rect 6620 3716 6628 3724
rect 6668 3716 6676 3724
rect 6716 3716 6724 3724
rect 6732 3716 6740 3724
rect 6796 3716 6804 3724
rect 6828 3716 6836 3724
rect 6860 3716 6868 3724
rect 6876 3716 6884 3724
rect 6924 3716 6932 3724
rect 6956 3716 6964 3724
rect 6972 3716 6980 3724
rect 7020 3716 7028 3724
rect 7052 3716 7060 3724
rect 7132 3716 7140 3724
rect 7196 3716 7204 3724
rect 7276 3716 7284 3724
rect 7324 3716 7332 3724
rect 7372 3716 7380 3724
rect 5740 3696 5748 3704
rect 6012 3696 6020 3704
rect 6124 3696 6132 3704
rect 6620 3696 6628 3704
rect 6652 3696 6660 3704
rect 6764 3696 6772 3704
rect 7164 3696 7172 3704
rect 7228 3696 7236 3704
rect 1276 3676 1284 3684
rect 1324 3676 1332 3684
rect 1388 3676 1396 3684
rect 1500 3676 1508 3684
rect 1564 3676 1572 3684
rect 1628 3676 1636 3684
rect 1804 3676 1812 3684
rect 1868 3676 1876 3684
rect 2076 3676 2084 3684
rect 2524 3676 2532 3684
rect 3068 3676 3076 3684
rect 3436 3676 3444 3684
rect 3580 3676 3588 3684
rect 3452 3656 3460 3664
rect 3612 3676 3620 3684
rect 3948 3676 3956 3684
rect 3964 3676 3972 3684
rect 4076 3676 4084 3684
rect 5324 3676 5332 3684
rect 5356 3676 5364 3684
rect 6156 3676 6164 3684
rect 7100 3676 7108 3684
rect 6796 3656 6804 3664
rect 7068 3656 7076 3664
rect 28 3636 36 3644
rect 204 3636 212 3644
rect 348 3636 356 3644
rect 588 3636 596 3644
rect 668 3636 676 3644
rect 732 3636 740 3644
rect 796 3636 804 3644
rect 1132 3636 1140 3644
rect 1228 3636 1236 3644
rect 1308 3636 1316 3644
rect 1468 3636 1476 3644
rect 1516 3636 1524 3644
rect 1580 3636 1588 3644
rect 1644 3636 1652 3644
rect 1820 3636 1828 3644
rect 1852 3636 1860 3644
rect 2140 3636 2148 3644
rect 2300 3636 2308 3644
rect 2588 3636 2596 3644
rect 2684 3636 2692 3644
rect 2748 3636 2756 3644
rect 4092 3636 4100 3644
rect 4204 3636 4212 3644
rect 6220 3636 6228 3644
rect 6988 3636 6996 3644
rect 7132 3636 7140 3644
rect 7244 3636 7252 3644
rect 7292 3636 7300 3644
rect 1411 3606 1419 3614
rect 1421 3606 1429 3614
rect 1431 3606 1439 3614
rect 1441 3606 1449 3614
rect 1451 3606 1459 3614
rect 1461 3606 1469 3614
rect 4419 3606 4427 3614
rect 4429 3606 4437 3614
rect 4439 3606 4447 3614
rect 4449 3606 4457 3614
rect 4459 3606 4467 3614
rect 4469 3606 4477 3614
rect 1052 3576 1060 3584
rect 1292 3576 1300 3584
rect 3036 3576 3044 3584
rect 3180 3576 3188 3584
rect 3388 3576 3396 3584
rect 3484 3576 3492 3584
rect 4140 3576 4148 3584
rect 4892 3576 4900 3584
rect 4988 3576 4996 3584
rect 5372 3576 5380 3584
rect 5852 3576 5860 3584
rect 6012 3576 6020 3584
rect 6716 3576 6724 3584
rect 3820 3556 3828 3564
rect 6348 3556 6356 3564
rect 6924 3556 6932 3564
rect 1116 3536 1124 3544
rect 1228 3536 1236 3544
rect 1324 3536 1332 3544
rect 1404 3536 1412 3544
rect 1548 3536 1556 3544
rect 1580 3536 1588 3544
rect 1772 3536 1780 3544
rect 1804 3536 1812 3544
rect 2364 3536 2372 3544
rect 4092 3536 4100 3544
rect 508 3516 516 3524
rect 700 3516 708 3524
rect 60 3496 68 3504
rect 92 3496 100 3504
rect 172 3496 180 3504
rect 220 3496 228 3504
rect 284 3496 292 3504
rect 316 3496 324 3504
rect 412 3496 420 3504
rect 460 3496 468 3504
rect 652 3496 660 3504
rect 76 3476 84 3484
rect 108 3476 116 3484
rect 220 3476 228 3484
rect 428 3476 436 3484
rect 540 3476 548 3484
rect 572 3476 580 3484
rect 748 3516 756 3524
rect 812 3516 820 3524
rect 1020 3516 1028 3524
rect 1084 3516 1092 3524
rect 1164 3516 1172 3524
rect 1180 3516 1188 3524
rect 1196 3516 1204 3524
rect 1340 3516 1348 3524
rect 1372 3516 1380 3524
rect 1612 3516 1620 3524
rect 1628 3516 1636 3524
rect 1708 3516 1716 3524
rect 1884 3516 1892 3524
rect 2076 3516 2084 3524
rect 2172 3516 2180 3524
rect 2300 3516 2308 3524
rect 2460 3516 2468 3524
rect 3100 3516 3108 3524
rect 3420 3516 3428 3524
rect 3788 3516 3796 3524
rect 3852 3516 3860 3524
rect 3868 3516 3876 3524
rect 3996 3516 4004 3524
rect 4076 3516 4084 3524
rect 4092 3516 4100 3524
rect 764 3496 772 3504
rect 892 3496 900 3504
rect 924 3496 932 3504
rect 972 3496 980 3504
rect 1004 3496 1012 3504
rect 1052 3496 1060 3504
rect 1100 3496 1108 3504
rect 1212 3496 1220 3504
rect 1260 3496 1268 3504
rect 1340 3496 1348 3504
rect 1388 3496 1396 3504
rect 1484 3496 1492 3504
rect 1516 3496 1524 3504
rect 1596 3496 1604 3504
rect 1628 3496 1636 3504
rect 1740 3496 1748 3504
rect 1820 3496 1828 3504
rect 1916 3496 1924 3504
rect 1948 3496 1956 3504
rect 2044 3496 2052 3504
rect 2076 3496 2084 3504
rect 2108 3496 2116 3504
rect 2252 3496 2260 3504
rect 2364 3496 2372 3504
rect 2396 3496 2404 3504
rect 2732 3496 2740 3504
rect 748 3476 756 3484
rect 844 3476 852 3484
rect 908 3476 916 3484
rect 1068 3476 1076 3484
rect 1148 3476 1156 3484
rect 1500 3476 1508 3484
rect 1660 3476 1668 3484
rect 1676 3476 1684 3484
rect 1724 3476 1732 3484
rect 1900 3476 1908 3484
rect 2060 3476 2068 3484
rect 2220 3476 2228 3484
rect 2332 3476 2340 3484
rect 2348 3476 2356 3484
rect 2492 3476 2500 3484
rect 2572 3476 2580 3484
rect 2620 3476 2628 3484
rect 2732 3476 2740 3484
rect 3132 3496 3140 3504
rect 3308 3496 3316 3504
rect 3436 3496 3444 3504
rect 3468 3496 3476 3504
rect 3564 3496 3572 3504
rect 3596 3496 3604 3504
rect 3676 3496 3684 3504
rect 3740 3496 3748 3504
rect 3916 3496 3924 3504
rect 3980 3496 3988 3504
rect 4124 3536 4132 3544
rect 4172 3536 4180 3544
rect 4812 3536 4820 3544
rect 5132 3536 5140 3544
rect 6364 3536 6372 3544
rect 6412 3536 6420 3544
rect 7180 3536 7188 3544
rect 4204 3516 4212 3524
rect 4220 3516 4228 3524
rect 4764 3516 4772 3524
rect 4124 3496 4132 3504
rect 4172 3496 4180 3504
rect 4476 3496 4484 3504
rect 6636 3516 6644 3524
rect 4668 3494 4676 3502
rect 4812 3496 4820 3504
rect 4844 3496 4852 3504
rect 4860 3496 4868 3504
rect 4924 3496 4932 3504
rect 5004 3496 5012 3504
rect 5020 3496 5028 3504
rect 5036 3496 5044 3504
rect 5100 3496 5108 3504
rect 5116 3496 5124 3504
rect 5212 3496 5220 3504
rect 5260 3494 5268 3502
rect 5340 3496 5348 3504
rect 5388 3496 5396 3504
rect 5404 3496 5412 3504
rect 5420 3496 5428 3504
rect 5516 3496 5524 3504
rect 5532 3496 5540 3504
rect 5628 3496 5636 3504
rect 5676 3496 5684 3504
rect 5692 3496 5700 3504
rect 5756 3496 5764 3504
rect 5804 3496 5812 3504
rect 5820 3496 5828 3504
rect 5900 3496 5908 3504
rect 6028 3496 6036 3504
rect 6044 3496 6052 3504
rect 6060 3496 6068 3504
rect 6108 3496 6116 3504
rect 6156 3496 6164 3504
rect 6220 3494 6228 3502
rect 6284 3496 6292 3504
rect 6396 3496 6404 3504
rect 6860 3516 6868 3524
rect 6540 3494 6548 3502
rect 6684 3496 6692 3504
rect 6748 3496 6756 3504
rect 6812 3496 6820 3504
rect 6908 3496 6916 3504
rect 7020 3496 7028 3504
rect 7116 3496 7124 3504
rect 7164 3496 7172 3504
rect 7292 3496 7300 3504
rect 2844 3476 2852 3484
rect 2860 3476 2868 3484
rect 3020 3476 3028 3484
rect 3068 3480 3076 3488
rect 3148 3476 3156 3484
rect 3244 3476 3252 3484
rect 12 3456 20 3464
rect 124 3456 132 3464
rect 236 3456 244 3464
rect 364 3456 372 3464
rect 556 3456 564 3464
rect 620 3456 628 3464
rect 684 3456 692 3464
rect 860 3456 868 3464
rect 972 3456 980 3464
rect 1116 3456 1124 3464
rect 1340 3456 1348 3464
rect 1948 3456 1956 3464
rect 1996 3456 2004 3464
rect 2012 3456 2020 3464
rect 2156 3456 2164 3464
rect 2220 3456 2228 3464
rect 172 3436 180 3444
rect 284 3436 292 3444
rect 380 3436 388 3444
rect 492 3436 500 3444
rect 508 3436 516 3444
rect 540 3436 548 3444
rect 604 3436 612 3444
rect 636 3436 644 3444
rect 668 3436 676 3444
rect 716 3436 724 3444
rect 796 3436 804 3444
rect 812 3436 820 3444
rect 876 3436 884 3444
rect 988 3436 996 3444
rect 1148 3436 1156 3444
rect 1212 3436 1220 3444
rect 1596 3436 1604 3444
rect 1660 3436 1668 3444
rect 1692 3436 1700 3444
rect 1820 3436 1828 3444
rect 2028 3436 2036 3444
rect 2172 3436 2180 3444
rect 2236 3436 2244 3444
rect 2444 3456 2452 3464
rect 2508 3456 2516 3464
rect 2588 3456 2596 3464
rect 2620 3456 2628 3464
rect 3292 3476 3300 3484
rect 3324 3476 3332 3484
rect 3356 3476 3364 3484
rect 3468 3476 3476 3484
rect 3644 3476 3652 3484
rect 3708 3480 3716 3488
rect 3724 3476 3732 3484
rect 3740 3476 3748 3484
rect 3804 3476 3812 3484
rect 3900 3476 3908 3484
rect 3932 3476 3940 3484
rect 3996 3476 4004 3484
rect 4044 3476 4052 3484
rect 4156 3476 4164 3484
rect 4252 3476 4260 3484
rect 4396 3476 4404 3484
rect 4492 3476 4500 3484
rect 4700 3476 4708 3484
rect 4732 3476 4740 3484
rect 4828 3476 4836 3484
rect 5052 3476 5060 3484
rect 5436 3476 5444 3484
rect 3372 3456 3380 3464
rect 3404 3456 3412 3464
rect 3548 3456 3556 3464
rect 3932 3456 3940 3464
rect 4284 3456 4292 3464
rect 4524 3456 4532 3464
rect 5484 3456 5492 3464
rect 5564 3456 5572 3464
rect 5612 3476 5620 3484
rect 5644 3476 5652 3484
rect 5708 3476 5716 3484
rect 5788 3456 5796 3464
rect 6092 3456 6100 3464
rect 6140 3476 6148 3484
rect 6572 3476 6580 3484
rect 6604 3476 6612 3484
rect 6652 3476 6660 3484
rect 6700 3476 6708 3484
rect 6764 3456 6772 3464
rect 6844 3456 6852 3464
rect 6892 3476 6900 3484
rect 7132 3476 7140 3484
rect 7276 3476 7284 3484
rect 7052 3456 7060 3464
rect 7164 3456 7172 3464
rect 2284 3436 2292 3444
rect 2316 3436 2324 3444
rect 2460 3436 2468 3444
rect 2604 3436 2612 3444
rect 2700 3436 2708 3444
rect 2812 3436 2820 3444
rect 2892 3436 2900 3444
rect 3868 3436 3876 3444
rect 4012 3436 4020 3444
rect 4076 3436 4084 3444
rect 4236 3436 4244 3444
rect 4508 3436 4516 3444
rect 4540 3436 4548 3444
rect 5452 3436 5460 3444
rect 5596 3436 5604 3444
rect 5724 3436 5732 3444
rect 6780 3436 6788 3444
rect 124 3416 132 3424
rect 236 3416 244 3424
rect 1996 3416 2004 3424
rect 2156 3416 2164 3424
rect 2444 3416 2452 3424
rect 2620 3416 2628 3424
rect 2915 3406 2923 3414
rect 2925 3406 2933 3414
rect 2935 3406 2943 3414
rect 2945 3406 2953 3414
rect 2955 3406 2963 3414
rect 2965 3406 2973 3414
rect 5923 3406 5931 3414
rect 5933 3406 5941 3414
rect 5943 3406 5951 3414
rect 5953 3406 5961 3414
rect 5963 3406 5971 3414
rect 5973 3406 5981 3414
rect 12 3396 20 3404
rect 2236 3396 2244 3404
rect 3068 3396 3076 3404
rect 12 3356 20 3364
rect 44 3356 52 3364
rect 76 3356 84 3364
rect 300 3356 308 3364
rect 524 3356 532 3364
rect 924 3376 932 3384
rect 1228 3376 1236 3384
rect 1452 3376 1460 3384
rect 1628 3376 1636 3384
rect 1692 3376 1700 3384
rect 620 3356 628 3364
rect 844 3356 852 3364
rect 1708 3356 1716 3364
rect 1884 3356 1892 3364
rect 1932 3356 1940 3364
rect 2188 3356 2196 3364
rect 2236 3356 2244 3364
rect 2252 3356 2260 3364
rect 2572 3356 2580 3364
rect 2972 3376 2980 3384
rect 3276 3376 3284 3384
rect 3484 3376 3492 3384
rect 3612 3376 3620 3384
rect 3900 3376 3908 3384
rect 3932 3376 3940 3384
rect 3996 3376 4004 3384
rect 4300 3376 4308 3384
rect 4364 3376 4372 3384
rect 4556 3376 4564 3384
rect 4764 3376 4772 3384
rect 4956 3376 4964 3384
rect 5372 3376 5380 3384
rect 5692 3376 5700 3384
rect 5916 3376 5924 3384
rect 5996 3376 6004 3384
rect 6188 3376 6196 3384
rect 6444 3376 6452 3384
rect 6524 3376 6532 3384
rect 6844 3376 6852 3384
rect 7180 3376 7188 3384
rect 7212 3376 7220 3384
rect 2716 3356 2724 3364
rect 2860 3356 2868 3364
rect 3068 3356 3076 3364
rect 3340 3356 3348 3364
rect 3532 3356 3540 3364
rect 3644 3356 3652 3364
rect 3708 3356 3716 3364
rect 4060 3356 4068 3364
rect 4172 3356 4180 3364
rect 4572 3356 4580 3364
rect 5084 3356 5092 3364
rect 6380 3356 6388 3364
rect 6780 3356 6788 3364
rect 7196 3356 7204 3364
rect 44 3336 52 3344
rect 124 3336 132 3344
rect 268 3336 276 3344
rect 668 3336 676 3344
rect 764 3336 772 3344
rect 972 3336 980 3344
rect 1260 3332 1268 3340
rect 1276 3336 1284 3344
rect 1516 3336 1524 3344
rect 1532 3336 1540 3344
rect 1692 3336 1700 3344
rect 2236 3336 2244 3344
rect 2284 3336 2292 3344
rect 2348 3336 2356 3344
rect 2588 3336 2596 3344
rect 2620 3336 2628 3344
rect 2700 3336 2708 3344
rect 2764 3336 2772 3344
rect 2940 3336 2948 3344
rect 3036 3336 3044 3344
rect 3244 3336 3252 3344
rect 3516 3336 3524 3344
rect 3548 3336 3556 3344
rect 3564 3336 3572 3344
rect 3676 3336 3684 3344
rect 3740 3336 3748 3344
rect 3932 3336 3940 3344
rect 3964 3336 3972 3344
rect 4044 3336 4052 3344
rect 4108 3336 4116 3344
rect 4204 3336 4212 3344
rect 4348 3336 4356 3344
rect 4412 3336 4420 3344
rect 4604 3336 4612 3344
rect 4796 3336 4804 3344
rect 4972 3336 4980 3344
rect 5068 3336 5076 3344
rect 5164 3336 5172 3344
rect 5212 3336 5220 3344
rect 5404 3336 5412 3344
rect 5468 3336 5476 3344
rect 5580 3336 5588 3344
rect 5676 3336 5684 3344
rect 5756 3336 5764 3344
rect 6156 3336 6164 3344
rect 6284 3336 6292 3344
rect 6348 3336 6356 3344
rect 6460 3336 6468 3344
rect 6812 3336 6820 3344
rect 7036 3336 7044 3344
rect 7100 3336 7108 3344
rect 7132 3336 7140 3344
rect 7164 3336 7172 3344
rect 76 3316 84 3324
rect 108 3316 116 3324
rect 140 3316 148 3324
rect 172 3316 180 3324
rect 332 3316 340 3324
rect 380 3316 388 3324
rect 412 3316 420 3324
rect 476 3316 484 3324
rect 556 3316 564 3324
rect 620 3316 628 3324
rect 668 3316 676 3324
rect 716 3316 724 3324
rect 780 3316 788 3324
rect 812 3316 820 3324
rect 844 3316 852 3324
rect 876 3316 884 3324
rect 956 3316 964 3324
rect 1004 3316 1012 3324
rect 1068 3316 1076 3324
rect 1132 3316 1140 3324
rect 1212 3316 1220 3324
rect 1308 3316 1316 3324
rect 1356 3316 1364 3324
rect 1500 3316 1508 3324
rect 1548 3316 1556 3324
rect 1628 3316 1636 3324
rect 1660 3316 1668 3324
rect 1788 3316 1796 3324
rect 1852 3316 1860 3324
rect 1932 3316 1940 3324
rect 1964 3316 1972 3324
rect 2012 3316 2020 3324
rect 2076 3316 2084 3324
rect 2156 3316 2164 3324
rect 2188 3316 2196 3324
rect 2284 3316 2292 3324
rect 2316 3316 2324 3324
rect 140 3296 148 3304
rect 460 3296 468 3304
rect 732 3296 740 3304
rect 796 3296 804 3304
rect 860 3296 868 3304
rect 988 3296 996 3304
rect 1052 3296 1060 3304
rect 1116 3296 1124 3304
rect 1292 3296 1300 3304
rect 1644 3296 1652 3304
rect 1660 3296 1668 3304
rect 1804 3296 1812 3304
rect 1868 3296 1876 3304
rect 2028 3296 2036 3304
rect 2092 3296 2100 3304
rect 2428 3316 2436 3324
rect 2508 3316 2516 3324
rect 2540 3316 2548 3324
rect 2556 3316 2564 3324
rect 2604 3316 2612 3324
rect 2636 3316 2644 3324
rect 2732 3316 2740 3324
rect 2812 3316 2820 3324
rect 3212 3318 3220 3326
rect 3308 3316 3316 3324
rect 3388 3316 3396 3324
rect 3452 3316 3460 3324
rect 3580 3316 3588 3324
rect 3612 3316 3620 3324
rect 3660 3316 3668 3324
rect 3708 3316 3716 3324
rect 3772 3318 3780 3326
rect 3836 3316 3844 3324
rect 3980 3316 3988 3324
rect 4028 3316 4036 3324
rect 4092 3316 4100 3324
rect 4156 3316 4164 3324
rect 4220 3316 4228 3324
rect 4332 3316 4340 3324
rect 4396 3316 4404 3324
rect 4524 3316 4532 3324
rect 4540 3316 4548 3324
rect 4636 3318 4644 3326
rect 4844 3316 4852 3324
rect 4892 3316 4900 3324
rect 4988 3316 4996 3324
rect 5004 3316 5012 3324
rect 2364 3296 2372 3304
rect 2412 3296 2420 3304
rect 2524 3296 2532 3304
rect 3404 3296 3412 3304
rect 3468 3296 3476 3304
rect 3484 3296 3492 3304
rect 3612 3296 3620 3304
rect 3996 3296 4004 3304
rect 4060 3296 4068 3304
rect 4284 3296 4292 3304
rect 4364 3296 4372 3304
rect 5116 3316 5124 3324
rect 5148 3316 5156 3324
rect 5180 3316 5188 3324
rect 5244 3318 5252 3326
rect 5452 3316 5460 3324
rect 5596 3316 5604 3324
rect 5612 3316 5620 3324
rect 5036 3296 5044 3304
rect 5724 3316 5732 3324
rect 5788 3318 5796 3326
rect 6092 3316 6100 3324
rect 6316 3318 6324 3326
rect 6412 3316 6420 3324
rect 6476 3316 6484 3324
rect 6492 3316 6500 3324
rect 6540 3316 6548 3324
rect 6652 3316 6660 3324
rect 6716 3318 6724 3326
rect 6796 3316 6804 3324
rect 6828 3316 6836 3324
rect 6908 3316 6916 3324
rect 6956 3316 6964 3324
rect 7036 3316 7044 3324
rect 5644 3296 5652 3304
rect 7148 3316 7156 3324
rect 7276 3316 7284 3324
rect 7308 3316 7316 3324
rect 7100 3296 7108 3304
rect 428 3276 436 3284
rect 476 3276 484 3284
rect 492 3276 500 3284
rect 700 3276 708 3284
rect 764 3276 772 3284
rect 860 3276 868 3284
rect 1020 3276 1028 3284
rect 1084 3276 1092 3284
rect 1148 3276 1156 3284
rect 1180 3276 1188 3284
rect 1324 3276 1332 3284
rect 1580 3276 1588 3284
rect 1612 3276 1620 3284
rect 1772 3276 1780 3284
rect 1836 3276 1844 3284
rect 1916 3276 1924 3284
rect 1996 3276 2004 3284
rect 2012 3276 2020 3284
rect 2060 3276 2068 3284
rect 2444 3276 2452 3284
rect 2492 3276 2500 3284
rect 3084 3276 3092 3284
rect 3372 3276 3380 3284
rect 3436 3276 3444 3284
rect 5564 3276 5572 3284
rect 5884 3276 5892 3284
rect 1468 3256 1476 3264
rect 1964 3256 1972 3264
rect 3388 3256 3396 3264
rect 3452 3256 3460 3264
rect 108 3236 116 3244
rect 476 3236 484 3244
rect 540 3236 548 3244
rect 716 3236 724 3244
rect 908 3236 916 3244
rect 1036 3236 1044 3244
rect 1100 3236 1108 3244
rect 1164 3236 1172 3244
rect 1340 3236 1348 3244
rect 1740 3236 1748 3244
rect 1852 3236 1860 3244
rect 1980 3236 1988 3244
rect 2460 3236 2468 3244
rect 2508 3236 2516 3244
rect 2828 3236 2836 3244
rect 3052 3236 3060 3244
rect 3532 3236 3540 3244
rect 4268 3236 4276 3244
rect 6524 3236 6532 3244
rect 6572 3236 6580 3244
rect 6588 3236 6596 3244
rect 6844 3236 6852 3244
rect 1411 3206 1419 3214
rect 1421 3206 1429 3214
rect 1431 3206 1439 3214
rect 1441 3206 1449 3214
rect 1451 3206 1459 3214
rect 1461 3206 1469 3214
rect 4419 3206 4427 3214
rect 4429 3206 4437 3214
rect 4439 3206 4447 3214
rect 4449 3206 4457 3214
rect 4459 3206 4467 3214
rect 4469 3206 4477 3214
rect 812 3176 820 3184
rect 876 3176 884 3184
rect 940 3176 948 3184
rect 1020 3176 1028 3184
rect 1372 3176 1380 3184
rect 1388 3176 1396 3184
rect 1516 3176 1524 3184
rect 1580 3176 1588 3184
rect 1644 3176 1652 3184
rect 1708 3176 1716 3184
rect 1836 3176 1844 3184
rect 1948 3176 1956 3184
rect 2012 3176 2020 3184
rect 2092 3176 2100 3184
rect 2140 3176 2148 3184
rect 2908 3176 2916 3184
rect 3420 3176 3428 3184
rect 3628 3176 3636 3184
rect 3804 3176 3812 3184
rect 4060 3176 4068 3184
rect 4284 3176 4292 3184
rect 4316 3176 4324 3184
rect 4684 3176 4692 3184
rect 4844 3176 4852 3184
rect 5644 3176 5652 3184
rect 5676 3176 5684 3184
rect 6444 3176 6452 3184
rect 6716 3176 6724 3184
rect 6956 3176 6964 3184
rect 6988 3176 6996 3184
rect 1244 3156 1252 3164
rect 2300 3156 2308 3164
rect 2380 3156 2388 3164
rect 2828 3156 2836 3164
rect 3740 3156 3748 3164
rect 4220 3156 4228 3164
rect 796 3136 804 3144
rect 876 3136 884 3144
rect 1148 3136 1156 3144
rect 1500 3136 1508 3144
rect 1596 3136 1604 3144
rect 1660 3136 1668 3144
rect 1724 3136 1732 3144
rect 1788 3136 1796 3144
rect 1820 3136 1828 3144
rect 1852 3136 1860 3144
rect 1948 3136 1956 3144
rect 1964 3136 1972 3144
rect 2108 3136 2116 3144
rect 2156 3136 2164 3144
rect 2220 3136 2228 3144
rect 2284 3136 2292 3144
rect 2444 3136 2452 3144
rect 2492 3136 2500 3144
rect 2556 3136 2564 3144
rect 2764 3136 2772 3144
rect 3404 3136 3412 3144
rect 3500 3136 3508 3144
rect 3644 3136 3652 3144
rect 3852 3136 3860 3144
rect 4204 3136 4212 3144
rect 4268 3136 4276 3144
rect 4492 3136 4500 3144
rect 5324 3136 5332 3144
rect 5452 3136 5460 3144
rect 6236 3136 6244 3144
rect 60 3096 68 3104
rect 108 3116 116 3124
rect 684 3116 692 3124
rect 748 3116 756 3124
rect 1116 3116 1124 3124
rect 1132 3116 1140 3124
rect 1324 3116 1332 3124
rect 2412 3116 2420 3124
rect 2524 3116 2532 3124
rect 2636 3116 2644 3124
rect 2780 3116 2788 3124
rect 2796 3116 2804 3124
rect 3532 3116 3540 3124
rect 3548 3116 3556 3124
rect 3612 3116 3620 3124
rect 3708 3116 3716 3124
rect 4156 3116 4164 3124
rect 4236 3116 4244 3124
rect 4300 3116 4308 3124
rect 5068 3116 5076 3124
rect 5132 3116 5140 3124
rect 5148 3116 5156 3124
rect 5228 3116 5236 3124
rect 5724 3116 5732 3124
rect 5756 3116 5764 3124
rect 204 3096 212 3104
rect 252 3096 260 3104
rect 268 3096 276 3104
rect 364 3096 372 3104
rect 396 3096 404 3104
rect 508 3096 516 3104
rect 556 3096 564 3104
rect 588 3096 596 3104
rect 700 3096 708 3104
rect 92 3076 100 3084
rect 140 3076 148 3084
rect 252 3076 260 3084
rect 652 3076 660 3084
rect 780 3076 788 3084
rect 812 3096 820 3104
rect 876 3096 884 3104
rect 924 3096 932 3104
rect 988 3096 996 3104
rect 1004 3096 1012 3104
rect 1068 3096 1076 3104
rect 1116 3096 1124 3104
rect 1148 3096 1156 3104
rect 1276 3096 1284 3104
rect 1340 3096 1348 3104
rect 1420 3096 1428 3104
rect 940 3076 948 3084
rect 1004 3076 1012 3084
rect 1020 3076 1028 3084
rect 1068 3076 1076 3084
rect 1196 3076 1204 3084
rect 1212 3080 1220 3088
rect 1260 3076 1268 3084
rect 1516 3096 1524 3104
rect 1580 3096 1588 3104
rect 1644 3096 1652 3104
rect 1708 3096 1716 3104
rect 1772 3096 1780 3104
rect 1836 3096 1844 3104
rect 1884 3096 1892 3104
rect 1948 3096 1956 3104
rect 1996 3096 2004 3104
rect 2060 3096 2068 3104
rect 2012 3076 2020 3084
rect 2092 3096 2100 3104
rect 2172 3096 2180 3104
rect 2236 3096 2244 3104
rect 2300 3096 2308 3104
rect 2332 3096 2340 3104
rect 2380 3076 2388 3084
rect 2428 3096 2436 3104
rect 2540 3096 2548 3104
rect 2668 3096 2676 3104
rect 2764 3096 2772 3104
rect 2828 3096 2836 3104
rect 2876 3096 2884 3104
rect 3020 3096 3028 3104
rect 3052 3096 3060 3104
rect 3292 3096 3300 3104
rect 3516 3096 3524 3104
rect 3548 3096 3556 3104
rect 3580 3096 3588 3104
rect 3628 3096 3636 3104
rect 3676 3096 3684 3104
rect 3724 3096 3732 3104
rect 3788 3096 3796 3104
rect 3948 3096 3956 3104
rect 3996 3094 4004 3102
rect 4156 3096 4164 3104
rect 4220 3096 4228 3104
rect 4284 3096 4292 3104
rect 4316 3096 4324 3104
rect 4364 3096 4372 3104
rect 4476 3096 4484 3104
rect 4588 3096 4596 3104
rect 4716 3096 4724 3104
rect 4780 3096 4788 3104
rect 4940 3096 4948 3104
rect 5068 3096 5076 3104
rect 5180 3096 5188 3104
rect 5196 3096 5204 3104
rect 5292 3096 5300 3104
rect 5340 3096 5348 3104
rect 5356 3096 5364 3104
rect 5388 3096 5396 3104
rect 5436 3096 5444 3104
rect 5452 3096 5460 3104
rect 5516 3096 5524 3104
rect 5612 3096 5620 3104
rect 5708 3096 5716 3104
rect 5772 3096 5780 3104
rect 5916 3094 5924 3102
rect 6044 3096 6052 3104
rect 6076 3096 6084 3104
rect 6140 3096 6148 3104
rect 6188 3096 6196 3104
rect 6236 3096 6244 3104
rect 6252 3096 6260 3104
rect 6300 3096 6308 3104
rect 6540 3116 6548 3124
rect 6364 3096 6372 3104
rect 6476 3096 6484 3104
rect 6572 3096 6580 3104
rect 6876 3116 6884 3124
rect 6636 3096 6644 3104
rect 6700 3096 6708 3104
rect 6764 3096 6772 3104
rect 6780 3096 6788 3104
rect 6844 3096 6852 3104
rect 6860 3096 6868 3104
rect 6956 3096 6964 3104
rect 7036 3096 7044 3104
rect 7148 3096 7156 3104
rect 7244 3096 7252 3104
rect 7308 3096 7316 3104
rect 7340 3096 7348 3104
rect 2588 3076 2596 3084
rect 3004 3076 3012 3084
rect 3036 3076 3044 3084
rect 3116 3076 3124 3084
rect 3212 3076 3220 3084
rect 3244 3076 3252 3084
rect 3452 3076 3460 3084
rect 3596 3076 3604 3084
rect 3676 3076 3684 3084
rect 3740 3076 3748 3084
rect 3772 3076 3780 3084
rect 4172 3076 4180 3084
rect 4364 3076 4372 3084
rect 4380 3076 4388 3084
rect 4604 3076 4612 3084
rect 4732 3076 4740 3084
rect 4764 3076 4772 3084
rect 4860 3076 4868 3084
rect 4892 3076 4900 3084
rect 5116 3076 5124 3084
rect 5164 3076 5172 3084
rect 5372 3076 5380 3084
rect 5452 3076 5460 3084
rect 5500 3076 5508 3084
rect 5564 3076 5572 3084
rect 5612 3076 5620 3084
rect 5884 3076 5892 3084
rect 6124 3076 6132 3084
rect 6252 3076 6260 3084
rect 6284 3076 6292 3084
rect 6316 3076 6324 3084
rect 6332 3076 6340 3084
rect 6380 3076 6388 3084
rect 6428 3076 6436 3084
rect 6460 3076 6468 3084
rect 6524 3076 6532 3084
rect 6588 3076 6596 3084
rect 6604 3076 6612 3084
rect 6652 3076 6660 3084
rect 6748 3076 6756 3084
rect 6908 3076 6916 3084
rect 6972 3076 6980 3084
rect 7020 3076 7028 3084
rect 7180 3076 7188 3084
rect 7260 3076 7268 3084
rect 7292 3076 7300 3084
rect 7340 3076 7348 3084
rect 12 3056 20 3064
rect 156 3056 164 3064
rect 300 3056 308 3064
rect 316 3056 324 3064
rect 364 3056 372 3064
rect 444 3056 452 3064
rect 460 3056 468 3064
rect 140 3036 148 3044
rect 204 3036 212 3044
rect 284 3036 292 3044
rect 476 3036 484 3044
rect 556 3056 564 3064
rect 620 3056 628 3064
rect 732 3056 740 3064
rect 924 3056 932 3064
rect 1004 3056 1012 3064
rect 1996 3056 2004 3064
rect 2508 3056 2516 3064
rect 2588 3056 2596 3064
rect 2716 3056 2724 3064
rect 668 3036 676 3044
rect 716 3036 724 3044
rect 748 3036 756 3044
rect 1068 3036 1076 3044
rect 1148 3036 1156 3044
rect 2556 3036 2564 3044
rect 2764 3036 2772 3044
rect 2972 3056 2980 3064
rect 3084 3056 3092 3064
rect 3420 3056 3428 3064
rect 3820 3056 3828 3064
rect 3852 3056 3860 3064
rect 3900 3056 3908 3064
rect 4076 3056 4084 3064
rect 4092 3056 4100 3064
rect 4348 3056 4356 3064
rect 4412 3056 4420 3064
rect 4700 3056 4708 3064
rect 4812 3056 4820 3064
rect 5484 3056 5492 3064
rect 5580 3056 5588 3064
rect 6076 3056 6084 3064
rect 6092 3056 6100 3064
rect 6204 3056 6212 3064
rect 6508 3056 6516 3064
rect 6668 3056 6676 3064
rect 6988 3056 6996 3064
rect 7308 3056 7316 3064
rect 7356 3056 7364 3064
rect 7388 3056 7396 3064
rect 3148 3036 3156 3044
rect 3836 3036 3844 3044
rect 5052 3036 5060 3044
rect 5388 3036 5396 3044
rect 5516 3036 5524 3044
rect 5788 3036 5796 3044
rect 6060 3036 6068 3044
rect 6812 3036 6820 3044
rect 7052 3036 7060 3044
rect 7276 3036 7284 3044
rect 12 3016 20 3024
rect 156 3016 164 3024
rect 316 3016 324 3024
rect 444 3016 452 3024
rect 2716 3016 2724 3024
rect 3084 3016 3092 3024
rect 2915 3006 2923 3014
rect 2925 3006 2933 3014
rect 2935 3006 2943 3014
rect 2945 3006 2953 3014
rect 2955 3006 2963 3014
rect 2965 3006 2973 3014
rect 5923 3006 5931 3014
rect 5933 3006 5941 3014
rect 5943 3006 5951 3014
rect 5953 3006 5961 3014
rect 5963 3006 5971 3014
rect 5973 3006 5981 3014
rect 204 2996 212 3004
rect 956 2996 964 3004
rect 1084 2996 1092 3004
rect 2268 2996 2276 3004
rect 2380 2996 2388 3004
rect 2492 2996 2500 3004
rect 2620 2996 2628 3004
rect 3020 2996 3028 3004
rect 140 2976 148 2984
rect 524 2976 532 2984
rect 844 2976 852 2984
rect 876 2976 884 2984
rect 908 2976 916 2984
rect 1196 2976 1204 2984
rect 1260 2976 1268 2984
rect 1308 2976 1316 2984
rect 1324 2976 1332 2984
rect 1500 2976 1508 2984
rect 1516 2976 1524 2984
rect 1644 2976 1652 2984
rect 1852 2976 1860 2984
rect 1900 2976 1908 2984
rect 2028 2976 2036 2984
rect 2108 2976 2116 2984
rect 2396 2976 2404 2984
rect 2444 2976 2452 2984
rect 2476 2976 2484 2984
rect 2540 2976 2548 2984
rect 2636 2976 2644 2984
rect 2668 2976 2676 2984
rect 2716 2976 2724 2984
rect 3372 2976 3380 2984
rect 3436 2976 3444 2984
rect 3500 2976 3508 2984
rect 3692 2976 3700 2984
rect 3788 2976 3796 2984
rect 4140 2976 4148 2984
rect 4300 2976 4308 2984
rect 4396 2976 4404 2984
rect 4540 2976 4548 2984
rect 4572 2976 4580 2984
rect 4604 2976 4612 2984
rect 4876 2976 4884 2984
rect 5212 2976 5220 2984
rect 5260 2976 5268 2984
rect 5628 2976 5636 2984
rect 5852 2976 5860 2984
rect 6108 2976 6116 2984
rect 6300 2976 6308 2984
rect 6364 2976 6372 2984
rect 6620 2976 6628 2984
rect 6780 2976 6788 2984
rect 12 2956 20 2964
rect 188 2956 196 2964
rect 204 2956 212 2964
rect 412 2956 420 2964
rect 588 2956 596 2964
rect 604 2956 612 2964
rect 636 2956 644 2964
rect 892 2956 900 2964
rect 956 2956 964 2964
rect 1004 2956 1012 2964
rect 1084 2956 1092 2964
rect 1356 2956 1364 2964
rect 1756 2956 1764 2964
rect 92 2936 100 2944
rect 140 2936 148 2944
rect 268 2936 276 2944
rect 524 2936 532 2944
rect 572 2936 580 2944
rect 812 2936 820 2944
rect 844 2936 852 2944
rect 1132 2936 1140 2944
rect 1196 2936 1204 2944
rect 1228 2936 1236 2944
rect 60 2916 68 2924
rect 156 2916 164 2924
rect 204 2916 212 2924
rect 252 2916 260 2924
rect 284 2916 292 2924
rect 364 2916 372 2924
rect 444 2916 452 2924
rect 476 2916 484 2924
rect 524 2916 532 2924
rect 588 2916 596 2924
rect 604 2916 612 2924
rect 636 2916 644 2924
rect 684 2916 692 2924
rect 764 2916 772 2924
rect 108 2896 116 2904
rect 348 2896 356 2904
rect 460 2896 468 2904
rect 700 2896 708 2904
rect 860 2916 868 2924
rect 940 2916 948 2924
rect 1004 2916 1012 2924
rect 1052 2916 1060 2924
rect 1084 2916 1092 2924
rect 1148 2916 1156 2924
rect 1308 2936 1316 2944
rect 1564 2936 1572 2944
rect 1660 2936 1668 2944
rect 1708 2936 1716 2944
rect 1740 2936 1748 2944
rect 1868 2936 1876 2944
rect 2044 2956 2052 2964
rect 2124 2956 2132 2964
rect 2236 2956 2244 2964
rect 2268 2956 2276 2964
rect 2300 2956 2308 2964
rect 2380 2956 2388 2964
rect 2492 2956 2500 2964
rect 2620 2956 2628 2964
rect 2732 2956 2740 2964
rect 2748 2956 2756 2964
rect 2780 2956 2788 2964
rect 2812 2956 2820 2964
rect 2908 2956 2916 2964
rect 3020 2956 3028 2964
rect 3100 2956 3108 2964
rect 3132 2956 3140 2964
rect 3388 2956 3396 2964
rect 3404 2956 3412 2964
rect 3452 2956 3460 2964
rect 3468 2956 3476 2964
rect 3484 2956 3492 2964
rect 3772 2956 3780 2964
rect 3964 2956 3972 2964
rect 4156 2956 4164 2964
rect 4268 2956 4276 2964
rect 4364 2956 4372 2964
rect 4508 2956 4516 2964
rect 4588 2956 4596 2964
rect 4748 2956 4756 2964
rect 2028 2936 2036 2944
rect 2044 2936 2052 2944
rect 2108 2936 2116 2944
rect 2140 2936 2148 2944
rect 2428 2936 2436 2944
rect 2444 2936 2452 2944
rect 2636 2936 2644 2944
rect 2716 2936 2724 2944
rect 2860 2936 2868 2944
rect 2892 2936 2900 2944
rect 2940 2936 2948 2944
rect 3276 2936 3284 2944
rect 3356 2936 3364 2944
rect 3516 2936 3524 2944
rect 3660 2936 3668 2944
rect 3692 2936 3700 2944
rect 3756 2936 3764 2944
rect 3788 2936 3796 2944
rect 3980 2936 3988 2944
rect 4076 2936 4084 2944
rect 4124 2936 4132 2944
rect 4188 2936 4196 2944
rect 4220 2936 4228 2944
rect 4316 2936 4324 2944
rect 4412 2936 4420 2944
rect 4524 2936 4532 2944
rect 4684 2936 4692 2944
rect 4892 2936 4900 2944
rect 5020 2936 5028 2944
rect 5052 2936 5060 2944
rect 5244 2936 5252 2944
rect 5292 2956 5300 2964
rect 5868 2956 5876 2964
rect 7020 2956 7028 2964
rect 5340 2936 5348 2944
rect 5404 2936 5412 2944
rect 5436 2936 5444 2944
rect 5468 2936 5476 2944
rect 5644 2936 5652 2944
rect 5980 2936 5988 2944
rect 6076 2936 6084 2944
rect 6156 2936 6164 2944
rect 6412 2936 6420 2944
rect 6476 2936 6484 2944
rect 6972 2936 6980 2944
rect 7068 2936 7076 2944
rect 7164 2936 7172 2944
rect 1260 2916 1268 2924
rect 1388 2916 1396 2924
rect 1468 2916 1476 2924
rect 1548 2916 1556 2924
rect 1612 2916 1620 2924
rect 1676 2916 1684 2924
rect 1692 2916 1700 2924
rect 1756 2916 1764 2924
rect 1804 2916 1812 2924
rect 1948 2916 1956 2924
rect 1980 2916 1988 2924
rect 2044 2916 2052 2924
rect 2060 2916 2068 2924
rect 2124 2916 2132 2924
rect 2140 2916 2148 2924
rect 2300 2916 2308 2924
rect 2332 2916 2340 2924
rect 2540 2916 2548 2924
rect 2588 2916 2596 2924
rect 2764 2916 2772 2924
rect 2876 2916 2884 2924
rect 3068 2916 3076 2924
rect 3196 2916 3204 2924
rect 3244 2916 3252 2924
rect 3260 2916 3268 2924
rect 3356 2916 3364 2924
rect 3532 2916 3540 2924
rect 3564 2916 3572 2924
rect 3628 2916 3636 2924
rect 3644 2916 3652 2924
rect 3676 2916 3684 2924
rect 3740 2916 3748 2924
rect 3804 2916 3812 2924
rect 3900 2916 3908 2924
rect 3964 2916 3972 2924
rect 4012 2916 4020 2924
rect 4076 2916 4084 2924
rect 4108 2916 4116 2924
rect 4172 2916 4180 2924
rect 4236 2916 4244 2924
rect 4284 2916 4292 2924
rect 4316 2916 4324 2924
rect 4332 2916 4340 2924
rect 4428 2916 4436 2924
rect 4764 2916 4772 2924
rect 5100 2916 5108 2924
rect 5228 2916 5236 2924
rect 5324 2916 5332 2924
rect 5340 2916 5348 2924
rect 5500 2918 5508 2926
rect 812 2896 820 2904
rect 1100 2896 1108 2904
rect 1196 2896 1204 2904
rect 1340 2896 1348 2904
rect 1596 2896 1604 2904
rect 1820 2896 1828 2904
rect 1868 2896 1876 2904
rect 1964 2896 1972 2904
rect 2188 2896 2196 2904
rect 2396 2896 2404 2904
rect 2476 2896 2484 2904
rect 2668 2896 2676 2904
rect 2700 2896 2708 2904
rect 2844 2896 2852 2904
rect 3084 2896 3092 2904
rect 3212 2896 3220 2904
rect 3228 2896 3236 2904
rect 3548 2896 3556 2904
rect 3612 2896 3620 2904
rect 3884 2896 3892 2904
rect 3948 2896 3956 2904
rect 4028 2896 4036 2904
rect 4092 2896 4100 2904
rect 4188 2896 4196 2904
rect 4380 2896 4388 2904
rect 4604 2896 4612 2904
rect 4636 2896 4644 2904
rect 5820 2916 5828 2924
rect 5836 2916 5844 2924
rect 5884 2916 5892 2924
rect 6028 2916 6036 2924
rect 6060 2916 6068 2924
rect 6172 2916 6180 2924
rect 6220 2916 6228 2924
rect 6284 2916 6292 2924
rect 6332 2916 6340 2924
rect 6348 2916 6356 2924
rect 6396 2916 6404 2924
rect 6444 2916 6452 2924
rect 6460 2916 6468 2924
rect 6508 2916 6516 2924
rect 6556 2916 6564 2924
rect 6572 2916 6580 2924
rect 6604 2916 6612 2924
rect 6652 2916 6660 2924
rect 6668 2916 6676 2924
rect 6700 2916 6708 2924
rect 6844 2916 6852 2924
rect 6892 2916 6900 2924
rect 7052 2916 7060 2924
rect 7116 2916 7124 2924
rect 7244 2916 7252 2924
rect 7276 2916 7284 2924
rect 5404 2896 5412 2904
rect 5900 2896 5908 2904
rect 5932 2896 5940 2904
rect 6364 2896 6372 2904
rect 6428 2896 6436 2904
rect 7004 2896 7012 2904
rect 380 2876 388 2884
rect 428 2876 436 2884
rect 492 2876 500 2884
rect 572 2876 580 2884
rect 668 2876 676 2884
rect 1132 2876 1140 2884
rect 1276 2876 1284 2884
rect 1772 2876 1780 2884
rect 1788 2876 1796 2884
rect 1932 2876 1940 2884
rect 2812 2876 2820 2884
rect 3052 2876 3060 2884
rect 3180 2876 3188 2884
rect 3580 2876 3588 2884
rect 3916 2876 3924 2884
rect 3932 2876 3940 2884
rect 4060 2876 4068 2884
rect 6204 2876 6212 2884
rect 6252 2876 6260 2884
rect 6988 2876 6996 2884
rect 7020 2876 7028 2884
rect 3564 2856 3572 2864
rect 364 2836 372 2844
rect 508 2836 516 2844
rect 1740 2836 1748 2844
rect 1916 2836 1924 2844
rect 2204 2836 2212 2844
rect 2828 2836 2836 2844
rect 2940 2836 2948 2844
rect 3068 2836 3076 2844
rect 3116 2836 3124 2844
rect 3148 2836 3156 2844
rect 3196 2836 3204 2844
rect 5756 2836 5764 2844
rect 5788 2836 5796 2844
rect 6028 2836 6036 2844
rect 6108 2836 6116 2844
rect 6540 2836 6548 2844
rect 6716 2836 6724 2844
rect 7084 2836 7092 2844
rect 7180 2836 7188 2844
rect 1411 2806 1419 2814
rect 1421 2806 1429 2814
rect 1431 2806 1439 2814
rect 1441 2806 1449 2814
rect 1451 2806 1459 2814
rect 1461 2806 1469 2814
rect 4419 2806 4427 2814
rect 4429 2806 4437 2814
rect 4439 2806 4447 2814
rect 4449 2806 4457 2814
rect 4459 2806 4467 2814
rect 4469 2806 4477 2814
rect 460 2776 468 2784
rect 780 2776 788 2784
rect 892 2776 900 2784
rect 940 2776 948 2784
rect 1084 2776 1092 2784
rect 1116 2776 1124 2784
rect 1292 2776 1300 2784
rect 1372 2776 1380 2784
rect 1516 2776 1524 2784
rect 1724 2776 1732 2784
rect 2716 2776 2724 2784
rect 2780 2776 2788 2784
rect 4108 2776 4116 2784
rect 4348 2776 4356 2784
rect 4380 2776 4388 2784
rect 4492 2776 4500 2784
rect 4540 2776 4548 2784
rect 4620 2776 4628 2784
rect 4668 2776 4676 2784
rect 4908 2776 4916 2784
rect 5932 2776 5940 2784
rect 6092 2776 6100 2784
rect 396 2736 404 2744
rect 444 2736 452 2744
rect 860 2756 868 2764
rect 2652 2756 2660 2764
rect 3516 2756 3524 2764
rect 4044 2756 4052 2764
rect 4172 2756 4180 2764
rect 60 2696 68 2704
rect 108 2716 116 2724
rect 524 2736 532 2744
rect 588 2736 596 2744
rect 796 2736 804 2744
rect 972 2736 980 2744
rect 1500 2736 1508 2744
rect 1740 2736 1748 2744
rect 2668 2736 2676 2744
rect 2732 2736 2740 2744
rect 2860 2736 2868 2744
rect 3372 2736 3380 2744
rect 3900 2736 3908 2744
rect 4156 2736 4164 2744
rect 4332 2736 4340 2744
rect 4556 2736 4564 2744
rect 5772 2736 5780 2744
rect 6268 2736 6276 2744
rect 6684 2736 6692 2744
rect 6924 2736 6932 2744
rect 7004 2736 7012 2744
rect 556 2716 564 2724
rect 908 2716 916 2724
rect 972 2716 980 2724
rect 1020 2716 1028 2724
rect 1068 2716 1076 2724
rect 1244 2716 1252 2724
rect 1708 2716 1716 2724
rect 1772 2716 1780 2724
rect 1804 2716 1812 2724
rect 1964 2716 1972 2724
rect 2140 2716 2148 2724
rect 2220 2716 2228 2724
rect 2444 2716 2452 2724
rect 2460 2716 2468 2724
rect 2636 2716 2644 2724
rect 2700 2716 2708 2724
rect 2812 2716 2820 2724
rect 2828 2716 2836 2724
rect 2940 2716 2948 2724
rect 3340 2716 3348 2724
rect 3420 2716 3428 2724
rect 3500 2716 3508 2724
rect 3596 2716 3604 2724
rect 3692 2716 3700 2724
rect 3900 2716 3908 2724
rect 4188 2716 4196 2724
rect 4204 2716 4212 2724
rect 4364 2716 4372 2724
rect 4652 2716 4660 2724
rect 4732 2716 4740 2724
rect 5148 2716 5156 2724
rect 5180 2716 5188 2724
rect 6204 2716 6212 2724
rect 6316 2716 6324 2724
rect 6556 2716 6564 2724
rect 204 2696 212 2704
rect 236 2696 244 2704
rect 300 2696 308 2704
rect 348 2696 356 2704
rect 412 2696 420 2704
rect 460 2696 468 2704
rect 92 2676 100 2684
rect 140 2676 148 2684
rect 348 2676 356 2684
rect 396 2676 404 2684
rect 508 2696 516 2704
rect 572 2696 580 2704
rect 668 2696 676 2704
rect 700 2696 708 2704
rect 780 2696 788 2704
rect 828 2696 836 2704
rect 1004 2696 1012 2704
rect 1148 2696 1156 2704
rect 1196 2696 1204 2704
rect 1500 2696 1508 2704
rect 1548 2696 1556 2704
rect 1564 2696 1572 2704
rect 1644 2696 1652 2704
rect 1676 2696 1684 2704
rect 1708 2696 1716 2704
rect 1756 2696 1764 2704
rect 1788 2696 1796 2704
rect 1836 2696 1844 2704
rect 2012 2696 2020 2704
rect 2044 2696 2052 2704
rect 2284 2696 2292 2704
rect 2332 2696 2340 2704
rect 2556 2696 2564 2704
rect 2652 2696 2660 2704
rect 2716 2696 2724 2704
rect 2780 2696 2788 2704
rect 2860 2696 2868 2704
rect 2988 2696 2996 2704
rect 3100 2696 3108 2704
rect 3260 2696 3268 2704
rect 3324 2696 3332 2704
rect 3356 2696 3364 2704
rect 3404 2696 3412 2704
rect 3468 2696 3476 2704
rect 3580 2696 3588 2704
rect 3836 2694 3844 2702
rect 3916 2696 3924 2704
rect 3964 2696 3972 2704
rect 4028 2696 4036 2704
rect 4092 2696 4100 2704
rect 4172 2696 4180 2704
rect 876 2676 884 2684
rect 924 2676 932 2684
rect 972 2676 980 2684
rect 1004 2676 1012 2684
rect 1164 2676 1172 2684
rect 1276 2676 1284 2684
rect 1436 2676 1444 2684
rect 1596 2680 1604 2688
rect 1612 2676 1620 2684
rect 1676 2676 1684 2684
rect 1868 2676 1876 2684
rect 2028 2676 2036 2684
rect 2108 2676 2116 2684
rect 2188 2676 2196 2684
rect 2412 2676 2420 2684
rect 2492 2676 2500 2684
rect 2540 2676 2548 2684
rect 2764 2676 2772 2684
rect 2876 2676 2884 2684
rect 3084 2676 3092 2684
rect 3212 2676 3220 2684
rect 3244 2676 3252 2684
rect 3260 2676 3268 2684
rect 3308 2676 3316 2684
rect 3356 2676 3364 2684
rect 3420 2676 3428 2684
rect 3452 2676 3460 2684
rect 3484 2676 3492 2684
rect 3596 2676 3604 2684
rect 3644 2676 3652 2684
rect 3660 2676 3668 2684
rect 4012 2676 4020 2684
rect 4076 2676 4084 2684
rect 4252 2696 4260 2704
rect 4268 2696 4276 2704
rect 4284 2696 4292 2704
rect 4348 2696 4356 2704
rect 4876 2696 4884 2704
rect 5004 2696 5012 2704
rect 5068 2694 5076 2702
rect 5148 2696 5156 2704
rect 5228 2696 5236 2704
rect 5372 2694 5380 2702
rect 5436 2696 5444 2704
rect 5484 2696 5492 2704
rect 5548 2696 5556 2704
rect 5644 2694 5652 2702
rect 5708 2696 5716 2704
rect 5804 2696 5812 2704
rect 5852 2696 5860 2704
rect 5868 2696 5876 2704
rect 5884 2696 5892 2704
rect 5900 2696 5908 2704
rect 6060 2696 6068 2704
rect 6108 2696 6116 2704
rect 6124 2696 6132 2704
rect 6140 2696 6148 2704
rect 6204 2696 6212 2704
rect 6252 2696 6260 2704
rect 6268 2696 6276 2704
rect 6364 2696 6372 2704
rect 6396 2696 6404 2704
rect 6428 2696 6436 2704
rect 6460 2696 6468 2704
rect 6524 2696 6532 2704
rect 6604 2716 6612 2724
rect 6668 2716 6676 2724
rect 6604 2696 6612 2704
rect 6796 2696 6804 2704
rect 6892 2696 6900 2704
rect 6972 2716 6980 2724
rect 7340 2716 7348 2724
rect 6972 2696 6980 2704
rect 7084 2696 7092 2704
rect 4300 2676 4308 2684
rect 4508 2676 4516 2684
rect 4588 2676 4596 2684
rect 4636 2676 4644 2684
rect 4684 2676 4692 2684
rect 4700 2676 4708 2684
rect 4748 2676 4756 2684
rect 4924 2676 4932 2684
rect 5132 2676 5140 2684
rect 5196 2676 5204 2684
rect 5404 2676 5412 2684
rect 5500 2676 5508 2684
rect 5548 2676 5556 2684
rect 6172 2676 6180 2684
rect 6188 2676 6196 2684
rect 6252 2676 6260 2684
rect 6364 2676 6372 2684
rect 6380 2676 6388 2684
rect 6444 2676 6452 2684
rect 6460 2676 6468 2684
rect 6508 2676 6516 2684
rect 6620 2676 6628 2684
rect 6636 2676 6644 2684
rect 6844 2676 6852 2684
rect 6876 2676 6884 2684
rect 6988 2676 6996 2684
rect 7116 2676 7124 2684
rect 7164 2676 7172 2684
rect 7196 2676 7204 2684
rect 7324 2676 7332 2684
rect 7372 2676 7380 2684
rect 12 2656 20 2664
rect 156 2656 164 2664
rect 236 2656 244 2664
rect 140 2636 148 2644
rect 332 2656 340 2664
rect 412 2656 420 2664
rect 620 2656 628 2664
rect 1180 2656 1188 2664
rect 1196 2656 1204 2664
rect 1308 2656 1316 2664
rect 1404 2656 1412 2664
rect 1628 2656 1636 2664
rect 1836 2656 1844 2664
rect 1852 2656 1860 2664
rect 1964 2656 1972 2664
rect 2092 2656 2100 2664
rect 2156 2656 2164 2664
rect 2236 2656 2244 2664
rect 2364 2656 2372 2664
rect 2396 2656 2404 2664
rect 2476 2656 2484 2664
rect 2524 2656 2532 2664
rect 3212 2656 3220 2664
rect 3276 2656 3284 2664
rect 3532 2656 3540 2664
rect 3548 2656 3556 2664
rect 3564 2656 3572 2664
rect 3836 2656 3844 2664
rect 3996 2656 4004 2664
rect 4012 2656 4020 2664
rect 4124 2656 4132 2664
rect 4460 2656 4468 2664
rect 4524 2656 4532 2664
rect 5468 2656 5476 2664
rect 5580 2656 5588 2664
rect 6300 2656 6308 2664
rect 6396 2656 6404 2664
rect 6492 2656 6500 2664
rect 316 2636 324 2644
rect 348 2636 356 2644
rect 604 2636 612 2644
rect 700 2636 708 2644
rect 860 2636 868 2644
rect 908 2636 916 2644
rect 1084 2636 1092 2644
rect 1244 2636 1252 2644
rect 1484 2636 1492 2644
rect 1916 2636 1924 2644
rect 2108 2636 2116 2644
rect 2140 2636 2148 2644
rect 2172 2636 2180 2644
rect 2188 2636 2196 2644
rect 2220 2636 2228 2644
rect 2284 2636 2292 2644
rect 2380 2636 2388 2644
rect 2412 2636 2420 2644
rect 2444 2636 2452 2644
rect 2540 2636 2548 2644
rect 3196 2636 3204 2644
rect 3676 2636 3684 2644
rect 3708 2636 3716 2644
rect 4572 2636 4580 2644
rect 4716 2636 4724 2644
rect 4940 2636 4948 2644
rect 5244 2636 5252 2644
rect 5452 2636 5460 2644
rect 5820 2636 5828 2644
rect 6316 2636 6324 2644
rect 6652 2636 6660 2644
rect 7340 2636 7348 2644
rect 620 2616 628 2624
rect 1964 2616 1972 2624
rect 2092 2616 2100 2624
rect 2156 2616 2164 2624
rect 2236 2616 2244 2624
rect 2364 2616 2372 2624
rect 2915 2606 2923 2614
rect 2925 2606 2933 2614
rect 2935 2606 2943 2614
rect 2945 2606 2953 2614
rect 2955 2606 2963 2614
rect 2965 2606 2973 2614
rect 5923 2606 5931 2614
rect 5933 2606 5941 2614
rect 5943 2606 5951 2614
rect 5953 2606 5961 2614
rect 5963 2606 5971 2614
rect 5973 2606 5981 2614
rect 12 2596 20 2604
rect 156 2596 164 2604
rect 988 2596 996 2604
rect 1100 2596 1108 2604
rect 1228 2596 1236 2604
rect 2412 2596 2420 2604
rect 2556 2596 2564 2604
rect 140 2576 148 2584
rect 620 2576 628 2584
rect 812 2576 820 2584
rect 1004 2576 1012 2584
rect 1340 2576 1348 2584
rect 1436 2576 1444 2584
rect 1500 2576 1508 2584
rect 1612 2576 1620 2584
rect 1692 2576 1700 2584
rect 1820 2576 1828 2584
rect 2204 2576 2212 2584
rect 2316 2576 2324 2584
rect 2636 2576 2644 2584
rect 2716 2576 2724 2584
rect 2828 2576 2836 2584
rect 3020 2576 3028 2584
rect 3644 2576 3652 2584
rect 3820 2576 3828 2584
rect 3948 2576 3956 2584
rect 4092 2576 4100 2584
rect 4540 2576 4548 2584
rect 4620 2576 4628 2584
rect 4764 2576 4772 2584
rect 4860 2576 4868 2584
rect 4892 2576 4900 2584
rect 4940 2576 4948 2584
rect 5180 2576 5188 2584
rect 5436 2576 5444 2584
rect 5868 2576 5876 2584
rect 6140 2576 6148 2584
rect 6412 2576 6420 2584
rect 6620 2576 6628 2584
rect 6988 2576 6996 2584
rect 7180 2576 7188 2584
rect 12 2556 20 2564
rect 156 2556 164 2564
rect 668 2556 676 2564
rect 988 2556 996 2564
rect 1084 2556 1092 2564
rect 1100 2556 1108 2564
rect 1228 2556 1236 2564
rect 1244 2556 1252 2564
rect 1420 2556 1428 2564
rect 1580 2556 1588 2564
rect 1628 2556 1636 2564
rect 1868 2556 1876 2564
rect 1932 2556 1940 2564
rect 2092 2556 2100 2564
rect 2252 2556 2260 2564
rect 2412 2556 2420 2564
rect 2428 2556 2436 2564
rect 2556 2556 2564 2564
rect 2812 2556 2820 2564
rect 2988 2556 2996 2564
rect 3116 2556 3124 2564
rect 3132 2556 3140 2564
rect 3564 2556 3572 2564
rect 3628 2556 3636 2564
rect 4012 2556 4020 2564
rect 4028 2556 4036 2564
rect 4044 2556 4052 2564
rect 4108 2556 4116 2564
rect 140 2536 148 2544
rect 60 2516 68 2524
rect 204 2516 212 2524
rect 220 2516 228 2524
rect 108 2496 116 2504
rect 316 2516 324 2524
rect 380 2516 388 2524
rect 460 2516 468 2524
rect 588 2536 596 2544
rect 620 2536 628 2544
rect 540 2516 548 2524
rect 252 2496 260 2504
rect 636 2516 644 2524
rect 716 2516 724 2524
rect 764 2516 772 2524
rect 828 2516 836 2524
rect 1164 2536 1172 2544
rect 1276 2536 1284 2544
rect 1516 2536 1524 2544
rect 1548 2536 1556 2544
rect 1740 2536 1748 2544
rect 1756 2536 1764 2544
rect 1852 2536 1860 2544
rect 1900 2536 1908 2544
rect 1948 2536 1956 2544
rect 1980 2536 1988 2544
rect 2012 2536 2020 2544
rect 2188 2536 2196 2544
rect 2236 2536 2244 2544
rect 2268 2536 2276 2544
rect 2316 2536 2324 2544
rect 2556 2536 2564 2544
rect 2668 2536 2676 2544
rect 2684 2536 2692 2544
rect 2780 2536 2788 2544
rect 2828 2536 2836 2544
rect 3100 2536 3108 2544
rect 3196 2536 3204 2544
rect 3596 2536 3604 2544
rect 3676 2536 3684 2544
rect 3724 2536 3732 2544
rect 3820 2536 3828 2544
rect 3868 2536 3876 2544
rect 3932 2536 3940 2544
rect 3980 2536 3988 2544
rect 4092 2536 4100 2544
rect 4140 2536 4148 2544
rect 4188 2536 4196 2544
rect 4220 2536 4228 2544
rect 4412 2536 4420 2544
rect 4700 2536 4708 2544
rect 4716 2536 4724 2544
rect 4780 2536 4788 2544
rect 4812 2536 4820 2544
rect 4828 2536 4836 2544
rect 4876 2536 4884 2544
rect 5004 2536 5012 2544
rect 5196 2536 5204 2544
rect 5212 2536 5220 2544
rect 5420 2536 5428 2544
rect 5468 2556 5476 2564
rect 5516 2556 5524 2564
rect 5532 2556 5540 2564
rect 5708 2556 5716 2564
rect 6060 2556 6068 2564
rect 5548 2536 5556 2544
rect 5852 2536 5860 2544
rect 6012 2536 6020 2544
rect 6332 2556 6340 2564
rect 7116 2556 7124 2564
rect 6108 2536 6116 2544
rect 6300 2536 6308 2544
rect 6364 2536 6372 2544
rect 6476 2536 6484 2544
rect 6540 2536 6548 2544
rect 6556 2536 6564 2544
rect 6860 2536 6868 2544
rect 6876 2536 6884 2544
rect 6972 2536 6980 2544
rect 588 2496 596 2504
rect 892 2496 900 2504
rect 924 2516 932 2524
rect 956 2516 964 2524
rect 1036 2516 1044 2524
rect 1052 2516 1060 2524
rect 1148 2516 1156 2524
rect 1180 2516 1188 2524
rect 1340 2516 1348 2524
rect 1388 2516 1396 2524
rect 1724 2516 1732 2524
rect 1900 2516 1908 2524
rect 1964 2516 1972 2524
rect 1996 2516 2004 2524
rect 2044 2516 2052 2524
rect 2172 2516 2180 2524
rect 2252 2516 2260 2524
rect 2316 2516 2324 2524
rect 2348 2516 2356 2524
rect 2364 2516 2372 2524
rect 2508 2516 2516 2524
rect 2844 2516 2852 2524
rect 3084 2516 3092 2524
rect 3260 2516 3268 2524
rect 3292 2516 3300 2524
rect 3436 2516 3444 2524
rect 3500 2518 3508 2526
rect 3564 2516 3572 2524
rect 3628 2516 3636 2524
rect 3660 2516 3668 2524
rect 3724 2516 3732 2524
rect 3756 2516 3764 2524
rect 3804 2516 3812 2524
rect 3868 2516 3876 2524
rect 3900 2516 3908 2524
rect 4156 2516 4164 2524
rect 4172 2516 4180 2524
rect 4236 2516 4244 2524
rect 4332 2516 4340 2524
rect 4508 2516 4516 2524
rect 4572 2516 4580 2524
rect 4732 2516 4740 2524
rect 5100 2516 5108 2524
rect 5228 2516 5236 2524
rect 5276 2516 5284 2524
rect 5308 2516 5316 2524
rect 5324 2516 5332 2524
rect 5372 2516 5380 2524
rect 5388 2516 5396 2524
rect 5404 2516 5412 2524
rect 5500 2516 5508 2524
rect 5564 2516 5572 2524
rect 5692 2516 5700 2524
rect 5804 2516 5812 2524
rect 5820 2516 5828 2524
rect 5900 2516 5908 2524
rect 5980 2516 5988 2524
rect 6028 2516 6036 2524
rect 6092 2516 6100 2524
rect 6124 2516 6132 2524
rect 6204 2516 6212 2524
rect 6252 2516 6260 2524
rect 6364 2516 6372 2524
rect 6380 2516 6388 2524
rect 6428 2516 6436 2524
rect 6492 2516 6500 2524
rect 6524 2516 6532 2524
rect 6588 2516 6596 2524
rect 6684 2516 6692 2524
rect 6732 2516 6740 2524
rect 6812 2516 6820 2524
rect 6844 2516 6852 2524
rect 1308 2496 1316 2504
rect 1516 2496 1524 2504
rect 1548 2496 1556 2504
rect 2028 2496 2036 2504
rect 2140 2496 2148 2504
rect 2204 2496 2212 2504
rect 2332 2496 2340 2504
rect 2476 2496 2484 2504
rect 3676 2496 3684 2504
rect 3756 2496 3764 2504
rect 3884 2496 3892 2504
rect 3948 2496 3956 2504
rect 3980 2496 3988 2504
rect 4092 2496 4100 2504
rect 4188 2496 4196 2504
rect 4604 2496 4612 2504
rect 4620 2496 4628 2504
rect 4652 2496 4660 2504
rect 4860 2496 4868 2504
rect 4908 2496 4916 2504
rect 4924 2496 4932 2504
rect 5100 2496 5108 2504
rect 5164 2496 5172 2504
rect 6492 2496 6500 2504
rect 6556 2496 6564 2504
rect 6812 2496 6820 2504
rect 6908 2496 6916 2504
rect 6956 2516 6964 2524
rect 7100 2516 7108 2524
rect 7244 2516 7252 2524
rect 7292 2516 7300 2524
rect 6956 2496 6964 2504
rect 332 2476 340 2484
rect 396 2476 404 2484
rect 444 2476 452 2484
rect 684 2476 692 2484
rect 780 2476 788 2484
rect 844 2476 852 2484
rect 988 2476 996 2484
rect 1244 2476 1252 2484
rect 1916 2476 1924 2484
rect 2060 2476 2068 2484
rect 3772 2476 3780 2484
rect 4252 2476 4260 2484
rect 4572 2476 4580 2484
rect 4604 2476 4612 2484
rect 4780 2476 4788 2484
rect 4956 2476 4964 2484
rect 5052 2476 5060 2484
rect 5340 2476 5348 2484
rect 5772 2456 5780 2464
rect 60 2436 68 2444
rect 316 2436 324 2444
rect 380 2436 388 2444
rect 460 2436 468 2444
rect 652 2436 660 2444
rect 764 2436 772 2444
rect 1068 2436 1076 2444
rect 1340 2436 1348 2444
rect 1676 2436 1684 2444
rect 2076 2436 2084 2444
rect 2124 2436 2132 2444
rect 2268 2436 2276 2444
rect 2460 2436 2468 2444
rect 3004 2436 3012 2444
rect 3164 2436 3172 2444
rect 3356 2436 3364 2444
rect 3372 2436 3380 2444
rect 3756 2436 3764 2444
rect 4540 2436 4548 2444
rect 5580 2436 5588 2444
rect 5868 2436 5876 2444
rect 6412 2436 6420 2444
rect 6460 2436 6468 2444
rect 7180 2436 7188 2444
rect 1411 2406 1419 2414
rect 1421 2406 1429 2414
rect 1431 2406 1439 2414
rect 1441 2406 1449 2414
rect 1451 2406 1459 2414
rect 1461 2406 1469 2414
rect 4419 2406 4427 2414
rect 4429 2406 4437 2414
rect 4439 2406 4447 2414
rect 4449 2406 4457 2414
rect 4459 2406 4467 2414
rect 4469 2406 4477 2414
rect 524 2376 532 2384
rect 1244 2376 1252 2384
rect 1564 2376 1572 2384
rect 1628 2376 1636 2384
rect 1900 2376 1908 2384
rect 2844 2376 2852 2384
rect 3020 2376 3028 2384
rect 3196 2376 3204 2384
rect 3628 2376 3636 2384
rect 3996 2376 4004 2384
rect 4092 2376 4100 2384
rect 4204 2376 4212 2384
rect 4524 2376 4532 2384
rect 4588 2376 4596 2384
rect 4668 2376 4676 2384
rect 6060 2376 6068 2384
rect 2044 2356 2052 2364
rect 3580 2356 3588 2364
rect 4636 2356 4644 2364
rect 380 2336 388 2344
rect 428 2336 436 2344
rect 572 2336 580 2344
rect 620 2336 628 2344
rect 780 2336 788 2344
rect 844 2336 852 2344
rect 876 2336 884 2344
rect 1004 2336 1012 2344
rect 1116 2336 1124 2344
rect 1548 2336 1556 2344
rect 1612 2336 1620 2344
rect 1692 2336 1700 2344
rect 2028 2336 2036 2344
rect 2156 2336 2164 2344
rect 2508 2336 2516 2344
rect 3276 2336 3284 2344
rect 3612 2336 3620 2344
rect 3980 2336 3988 2344
rect 3996 2336 4004 2344
rect 4124 2336 4132 2344
rect 4268 2336 4276 2344
rect 4396 2336 4404 2344
rect 4620 2336 4628 2344
rect 4716 2336 4724 2344
rect 5436 2336 5444 2344
rect 5804 2336 5812 2344
rect 6972 2336 6980 2344
rect 252 2316 260 2324
rect 364 2316 372 2324
rect 540 2316 548 2324
rect 1036 2316 1044 2324
rect 1420 2316 1428 2324
rect 1580 2316 1588 2324
rect 1644 2316 1652 2324
rect 1660 2316 1668 2324
rect 1964 2316 1972 2324
rect 2124 2316 2132 2324
rect 2268 2316 2276 2324
rect 2748 2316 2756 2324
rect 2780 2316 2788 2324
rect 2972 2316 2980 2324
rect 3052 2316 3060 2324
rect 3116 2316 3124 2324
rect 3228 2316 3236 2324
rect 3244 2316 3252 2324
rect 3532 2316 3540 2324
rect 3644 2316 3652 2324
rect 3708 2316 3716 2324
rect 3788 2316 3796 2324
rect 3852 2316 3860 2324
rect 4012 2316 4020 2324
rect 4268 2316 4276 2324
rect 4428 2316 4436 2324
rect 4652 2316 4660 2324
rect 4716 2316 4724 2324
rect 5084 2316 5092 2324
rect 5148 2316 5156 2324
rect 5500 2316 5508 2324
rect 5532 2316 5540 2324
rect 6284 2316 6292 2324
rect 6492 2316 6500 2324
rect 6524 2316 6532 2324
rect 44 2296 52 2304
rect 108 2296 116 2304
rect 140 2296 148 2304
rect 236 2296 244 2304
rect 284 2296 292 2304
rect 364 2296 372 2304
rect 412 2296 420 2304
rect 492 2296 500 2304
rect 524 2296 532 2304
rect 556 2296 564 2304
rect 604 2296 612 2304
rect 668 2296 676 2304
rect 716 2296 724 2304
rect 124 2276 132 2284
rect 428 2276 436 2284
rect 476 2276 484 2284
rect 572 2276 580 2284
rect 620 2276 628 2284
rect 668 2276 676 2284
rect 732 2276 740 2284
rect 764 2296 772 2304
rect 764 2276 772 2284
rect 828 2296 836 2304
rect 908 2296 916 2304
rect 956 2296 964 2304
rect 1020 2296 1028 2304
rect 1084 2296 1092 2304
rect 1132 2296 1140 2304
rect 1164 2296 1172 2304
rect 1228 2296 1236 2304
rect 1276 2296 1284 2304
rect 1308 2296 1316 2304
rect 1564 2296 1572 2304
rect 1628 2296 1636 2304
rect 1660 2296 1668 2304
rect 1740 2296 1748 2304
rect 1868 2296 1876 2304
rect 1900 2296 1908 2304
rect 2044 2296 2052 2304
rect 972 2276 980 2284
rect 1052 2276 1060 2284
rect 1180 2276 1188 2284
rect 12 2256 20 2264
rect 76 2256 84 2264
rect 188 2256 196 2264
rect 204 2256 212 2264
rect 412 2256 420 2264
rect 492 2256 500 2264
rect 604 2256 612 2264
rect 1100 2256 1108 2264
rect 1292 2276 1300 2284
rect 1340 2276 1348 2284
rect 1452 2276 1460 2284
rect 1692 2276 1700 2284
rect 1772 2276 1780 2284
rect 1996 2276 2004 2284
rect 2108 2296 2116 2304
rect 2140 2296 2148 2304
rect 2188 2296 2196 2304
rect 2268 2296 2276 2304
rect 2348 2296 2356 2304
rect 2396 2296 2404 2304
rect 2444 2296 2452 2304
rect 2540 2296 2548 2304
rect 2748 2296 2756 2304
rect 2780 2296 2788 2304
rect 3020 2296 3028 2304
rect 3084 2296 3092 2304
rect 3148 2296 3156 2304
rect 3276 2296 3284 2304
rect 3372 2296 3380 2304
rect 3436 2294 3444 2302
rect 3500 2296 3508 2304
rect 3548 2296 3556 2304
rect 3628 2296 3636 2304
rect 3676 2296 3684 2304
rect 3772 2296 3780 2304
rect 3804 2296 3812 2304
rect 3820 2296 3828 2304
rect 3916 2296 3924 2304
rect 3932 2296 3940 2304
rect 3996 2296 4004 2304
rect 4172 2296 4180 2304
rect 4316 2296 4324 2304
rect 4412 2296 4420 2304
rect 4556 2296 4564 2304
rect 4636 2296 4644 2304
rect 4700 2296 4708 2304
rect 4748 2296 4756 2304
rect 4796 2296 4804 2304
rect 4812 2296 4820 2304
rect 4956 2294 4964 2302
rect 5068 2296 5076 2304
rect 5084 2296 5092 2304
rect 5116 2296 5124 2304
rect 5180 2296 5188 2304
rect 5228 2296 5236 2304
rect 5276 2296 5284 2304
rect 5292 2296 5300 2304
rect 5324 2296 5332 2304
rect 5372 2296 5380 2304
rect 5388 2296 5396 2304
rect 5436 2296 5444 2304
rect 5452 2296 5460 2304
rect 5500 2296 5508 2304
rect 5564 2296 5572 2304
rect 5612 2296 5620 2304
rect 5660 2296 5668 2304
rect 5676 2296 5684 2304
rect 5724 2296 5732 2304
rect 5788 2296 5796 2304
rect 5868 2296 5876 2304
rect 5916 2296 5924 2304
rect 6092 2296 6100 2304
rect 6108 2296 6116 2304
rect 6172 2296 6180 2304
rect 6268 2296 6276 2304
rect 6284 2296 6292 2304
rect 6316 2296 6324 2304
rect 6364 2296 6372 2304
rect 6412 2296 6420 2304
rect 6460 2296 6468 2304
rect 6524 2296 6532 2304
rect 6556 2296 6564 2304
rect 6620 2296 6628 2304
rect 6636 2296 6644 2304
rect 6652 2296 6660 2304
rect 6700 2296 6708 2304
rect 6844 2296 6852 2304
rect 6940 2296 6948 2304
rect 7100 2296 7108 2304
rect 7244 2296 7252 2304
rect 7308 2294 7316 2302
rect 2140 2276 2148 2284
rect 2204 2276 2212 2284
rect 2252 2276 2260 2284
rect 2300 2276 2308 2284
rect 2348 2276 2356 2284
rect 2396 2276 2404 2284
rect 2428 2276 2436 2284
rect 2556 2276 2564 2284
rect 2572 2276 2580 2284
rect 2668 2276 2676 2284
rect 2700 2276 2708 2284
rect 2796 2276 2804 2284
rect 2812 2276 2820 2284
rect 2908 2276 2916 2284
rect 3036 2276 3044 2284
rect 3100 2276 3108 2284
rect 3164 2276 3172 2284
rect 3292 2276 3300 2284
rect 3420 2276 3428 2284
rect 3500 2276 3508 2284
rect 3660 2276 3668 2284
rect 3756 2276 3764 2284
rect 3836 2276 3844 2284
rect 3884 2276 3892 2284
rect 3948 2276 3956 2284
rect 4156 2276 4164 2284
rect 4396 2276 4404 2284
rect 4460 2276 4468 2284
rect 4748 2276 4756 2284
rect 4988 2276 4996 2284
rect 5052 2276 5060 2284
rect 5068 2276 5076 2284
rect 5132 2276 5140 2284
rect 5196 2276 5204 2284
rect 5212 2276 5220 2284
rect 5452 2276 5460 2284
rect 5516 2276 5524 2284
rect 5580 2276 5588 2284
rect 5756 2276 5764 2284
rect 5772 2276 5780 2284
rect 6028 2276 6036 2284
rect 6156 2276 6164 2284
rect 6188 2276 6196 2284
rect 6236 2276 6244 2284
rect 6332 2276 6340 2284
rect 6444 2276 6452 2284
rect 6572 2276 6580 2284
rect 6892 2276 6900 2284
rect 6924 2276 6932 2284
rect 7116 2276 7124 2284
rect 1212 2256 1220 2264
rect 1308 2256 1316 2264
rect 1340 2256 1348 2264
rect 1756 2256 1764 2264
rect 28 2236 36 2244
rect 380 2236 388 2244
rect 476 2236 484 2244
rect 668 2236 676 2244
rect 684 2236 692 2244
rect 828 2236 836 2244
rect 924 2236 932 2244
rect 1020 2236 1028 2244
rect 1692 2236 1700 2244
rect 2076 2256 2084 2264
rect 2108 2256 2116 2264
rect 2188 2256 2196 2264
rect 2316 2256 2324 2264
rect 2348 2256 2356 2264
rect 2380 2256 2388 2264
rect 2476 2256 2484 2264
rect 2684 2256 2692 2264
rect 4044 2256 4052 2264
rect 4076 2256 4084 2264
rect 4108 2256 4116 2264
rect 4204 2256 4212 2264
rect 4268 2256 4276 2264
rect 4300 2256 4308 2264
rect 4364 2256 4372 2264
rect 5020 2256 5028 2264
rect 5356 2256 5364 2264
rect 5404 2256 5412 2264
rect 5532 2256 5540 2264
rect 5692 2256 5700 2264
rect 6236 2256 6244 2264
rect 6380 2256 6388 2264
rect 6588 2256 6596 2264
rect 6668 2256 6676 2264
rect 1964 2236 1972 2244
rect 1996 2236 2004 2244
rect 2220 2236 2228 2244
rect 2252 2236 2260 2244
rect 2268 2236 2276 2244
rect 2604 2236 2612 2244
rect 3052 2236 3060 2244
rect 3116 2236 3124 2244
rect 3308 2236 3316 2244
rect 3740 2236 3748 2244
rect 4060 2236 4068 2244
rect 4124 2236 4132 2244
rect 4252 2236 4260 2244
rect 4828 2236 4836 2244
rect 5148 2236 5156 2244
rect 5628 2236 5636 2244
rect 6604 2236 6612 2244
rect 6732 2236 6740 2244
rect 6972 2236 6980 2244
rect 7180 2236 7188 2244
rect 76 2216 84 2224
rect 188 2216 196 2224
rect 204 2216 212 2224
rect 2316 2216 2324 2224
rect 2476 2216 2484 2224
rect 2915 2206 2923 2214
rect 2925 2206 2933 2214
rect 2935 2206 2943 2214
rect 2945 2206 2953 2214
rect 2955 2206 2963 2214
rect 2965 2206 2973 2214
rect 5923 2206 5931 2214
rect 5933 2206 5941 2214
rect 5943 2206 5951 2214
rect 5953 2206 5961 2214
rect 5963 2206 5971 2214
rect 5973 2206 5981 2214
rect 140 2176 148 2184
rect 332 2176 340 2184
rect 364 2176 372 2184
rect 460 2176 468 2184
rect 556 2176 564 2184
rect 588 2176 596 2184
rect 844 2176 852 2184
rect 1068 2176 1076 2184
rect 1212 2176 1220 2184
rect 1356 2176 1364 2184
rect 1916 2176 1924 2184
rect 2508 2176 2516 2184
rect 2540 2176 2548 2184
rect 2636 2176 2644 2184
rect 2748 2176 2756 2184
rect 2844 2176 2852 2184
rect 3068 2176 3076 2184
rect 3628 2176 3636 2184
rect 3676 2176 3684 2184
rect 3724 2176 3732 2184
rect 3788 2176 3796 2184
rect 3884 2176 3892 2184
rect 3932 2176 3940 2184
rect 4076 2176 4084 2184
rect 4108 2176 4116 2184
rect 4220 2176 4228 2184
rect 4284 2176 4292 2184
rect 4300 2176 4308 2184
rect 4460 2176 4468 2184
rect 4492 2176 4500 2184
rect 4556 2176 4564 2184
rect 4668 2176 4676 2184
rect 4764 2176 4772 2184
rect 5116 2176 5124 2184
rect 5468 2176 5476 2184
rect 5644 2176 5652 2184
rect 5868 2176 5876 2184
rect 5884 2176 5892 2184
rect 6044 2176 6052 2184
rect 6060 2176 6068 2184
rect 6172 2176 6180 2184
rect 6364 2176 6372 2184
rect 6924 2176 6932 2184
rect 76 2156 84 2164
rect 252 2156 260 2164
rect 268 2156 276 2164
rect 652 2156 660 2164
rect 1420 2156 1428 2164
rect 2092 2156 2100 2164
rect 2524 2156 2532 2164
rect 2684 2156 2692 2164
rect 2716 2156 2724 2164
rect 3404 2156 3412 2164
rect 3436 2156 3444 2164
rect 3468 2156 3476 2164
rect 3692 2156 3700 2164
rect 4476 2156 4484 2164
rect 4540 2156 4548 2164
rect 4636 2156 4644 2164
rect 5180 2156 5188 2164
rect 5612 2156 5620 2164
rect 92 2136 100 2144
rect 140 2136 148 2144
rect 172 2136 180 2144
rect 348 2136 356 2144
rect 364 2136 372 2144
rect 572 2136 580 2144
rect 588 2136 596 2144
rect 748 2136 756 2144
rect 892 2136 900 2144
rect 28 2116 36 2124
rect 76 2116 84 2124
rect 140 2116 148 2124
rect 188 2116 196 2124
rect 220 2116 228 2124
rect 252 2116 260 2124
rect 300 2116 308 2124
rect 396 2116 404 2124
rect 428 2116 436 2124
rect 476 2116 484 2124
rect 508 2116 516 2124
rect 620 2116 628 2124
rect 652 2116 660 2124
rect 732 2116 740 2124
rect 796 2116 804 2124
rect 812 2116 820 2124
rect 860 2116 868 2124
rect 940 2116 948 2124
rect 1004 2116 1012 2124
rect 1068 2116 1076 2124
rect 1132 2116 1140 2124
rect 1212 2136 1220 2144
rect 1356 2136 1364 2144
rect 1404 2136 1412 2144
rect 1196 2116 1204 2124
rect 1244 2116 1252 2124
rect 1308 2116 1316 2124
rect 1356 2116 1364 2124
rect 1420 2116 1428 2124
rect 1532 2116 1540 2124
rect 1628 2136 1636 2144
rect 1580 2116 1588 2124
rect 1644 2116 1652 2124
rect 1692 2116 1700 2124
rect 1724 2116 1732 2124
rect 1788 2116 1796 2124
rect 1996 2136 2004 2144
rect 1852 2116 1860 2124
rect 1916 2116 1924 2124
rect 1948 2116 1956 2124
rect 2252 2136 2260 2144
rect 2044 2116 2052 2124
rect 2156 2116 2164 2124
rect 2204 2116 2212 2124
rect 2332 2132 2340 2140
rect 2364 2136 2372 2144
rect 2460 2136 2468 2144
rect 2572 2136 2580 2144
rect 2668 2136 2676 2144
rect 2764 2136 2772 2144
rect 2780 2136 2788 2144
rect 2876 2136 2884 2144
rect 2956 2136 2964 2144
rect 3052 2136 3060 2144
rect 2556 2116 2564 2124
rect 2716 2116 2724 2124
rect 3116 2136 3124 2144
rect 3212 2136 3220 2144
rect 3228 2136 3236 2144
rect 3308 2136 3316 2144
rect 3372 2136 3380 2144
rect 3484 2136 3492 2144
rect 3580 2136 3588 2144
rect 3772 2136 3780 2144
rect 3836 2136 3844 2144
rect 3980 2136 3988 2144
rect 4092 2136 4100 2144
rect 4156 2136 4164 2144
rect 4188 2132 4196 2140
rect 4236 2136 4244 2144
rect 4348 2136 4356 2144
rect 4364 2136 4372 2144
rect 4588 2132 4596 2140
rect 4604 2136 4612 2144
rect 4652 2136 4660 2144
rect 4716 2136 4724 2144
rect 4732 2136 4740 2144
rect 4844 2136 4852 2144
rect 4972 2136 4980 2144
rect 5004 2136 5012 2144
rect 5068 2136 5076 2144
rect 5100 2136 5108 2144
rect 5484 2136 5492 2144
rect 5740 2156 5748 2164
rect 6380 2156 6388 2164
rect 6684 2156 6692 2164
rect 5660 2136 5668 2144
rect 5932 2136 5940 2144
rect 5980 2136 5988 2144
rect 6108 2136 6116 2144
rect 6124 2136 6132 2144
rect 6204 2136 6212 2144
rect 6412 2136 6420 2144
rect 6460 2136 6468 2144
rect 6524 2136 6532 2144
rect 6620 2136 6628 2144
rect 6716 2136 6724 2144
rect 6764 2136 6772 2144
rect 6796 2136 6804 2144
rect 6908 2136 6916 2144
rect 7084 2136 7092 2144
rect 12 2096 20 2104
rect 204 2096 212 2104
rect 316 2096 324 2104
rect 396 2096 404 2104
rect 412 2096 420 2104
rect 524 2096 532 2104
rect 540 2096 548 2104
rect 620 2096 628 2104
rect 636 2096 644 2104
rect 1244 2096 1252 2104
rect 1404 2096 1412 2104
rect 44 2076 52 2084
rect 92 2076 100 2084
rect 172 2076 180 2084
rect 444 2076 452 2084
rect 492 2076 500 2084
rect 668 2076 676 2084
rect 700 2076 708 2084
rect 924 2076 932 2084
rect 988 2076 996 2084
rect 1052 2076 1060 2084
rect 1116 2076 1124 2084
rect 1516 2076 1524 2084
rect 1868 2096 1876 2104
rect 1932 2096 1940 2104
rect 2028 2096 2036 2104
rect 2172 2096 2180 2104
rect 2188 2096 2196 2104
rect 2252 2096 2260 2104
rect 2508 2096 2516 2104
rect 2732 2096 2740 2104
rect 3260 2116 3268 2124
rect 3308 2116 3316 2124
rect 3516 2116 3524 2124
rect 3548 2116 3556 2124
rect 3644 2116 3652 2124
rect 3788 2116 3796 2124
rect 3916 2116 3924 2124
rect 3964 2116 3972 2124
rect 4028 2116 4036 2124
rect 4140 2116 4148 2124
rect 4252 2116 4260 2124
rect 4332 2116 4340 2124
rect 4700 2116 4708 2124
rect 4876 2116 4884 2124
rect 3276 2096 3284 2104
rect 3532 2096 3540 2104
rect 3628 2096 3636 2104
rect 3724 2096 3732 2104
rect 3788 2096 3796 2104
rect 3836 2096 3844 2104
rect 3868 2096 3876 2104
rect 3932 2096 3940 2104
rect 4044 2096 4052 2104
rect 4060 2096 4068 2104
rect 4396 2096 4404 2104
rect 4620 2096 4628 2104
rect 4764 2096 4772 2104
rect 5004 2096 5012 2104
rect 5052 2116 5060 2124
rect 5068 2116 5076 2124
rect 5148 2116 5156 2124
rect 5228 2116 5236 2124
rect 5244 2116 5252 2124
rect 5260 2116 5268 2124
rect 5324 2116 5332 2124
rect 5340 2116 5348 2124
rect 5356 2116 5364 2124
rect 5404 2116 5412 2124
rect 5436 2116 5444 2124
rect 5516 2116 5524 2124
rect 5564 2116 5572 2124
rect 5580 2116 5588 2124
rect 5676 2116 5684 2124
rect 5756 2116 5764 2124
rect 5916 2116 5924 2124
rect 6092 2116 6100 2124
rect 6140 2116 6148 2124
rect 6268 2116 6276 2124
rect 6428 2116 6436 2124
rect 6044 2096 6052 2104
rect 6460 2096 6468 2104
rect 6508 2116 6516 2124
rect 6572 2116 6580 2124
rect 6588 2116 6596 2124
rect 6636 2116 6644 2124
rect 6716 2116 6724 2124
rect 6780 2116 6788 2124
rect 6812 2116 6820 2124
rect 6844 2096 6852 2104
rect 6876 2116 6884 2124
rect 6892 2116 6900 2124
rect 7036 2116 7044 2124
rect 7148 2116 7156 2124
rect 7244 2116 7252 2124
rect 7260 2116 7268 2124
rect 1436 2056 1444 2064
rect 1596 2076 1604 2084
rect 1708 2076 1716 2084
rect 1772 2076 1780 2084
rect 1836 2076 1844 2084
rect 1900 2076 1908 2084
rect 2060 2076 2068 2084
rect 2140 2076 2148 2084
rect 2220 2076 2228 2084
rect 4012 2076 4020 2084
rect 4924 2076 4932 2084
rect 4972 2076 4980 2084
rect 6332 2076 6340 2084
rect 6428 2076 6436 2084
rect 7116 2076 7124 2084
rect 1676 2056 1684 2064
rect 1852 2056 1860 2064
rect 1996 2056 2004 2064
rect 4028 2056 4036 2064
rect 60 2036 68 2044
rect 236 2036 244 2044
rect 764 2036 772 2044
rect 908 2036 916 2044
rect 1004 2036 1012 2044
rect 1132 2036 1140 2044
rect 1228 2036 1236 2044
rect 1292 2036 1300 2044
rect 1340 2036 1348 2044
rect 1788 2036 1796 2044
rect 2076 2036 2084 2044
rect 2108 2036 2116 2044
rect 2156 2036 2164 2044
rect 2204 2036 2212 2044
rect 3420 2036 3428 2044
rect 3708 2036 3716 2044
rect 5196 2036 5204 2044
rect 5292 2036 5300 2044
rect 5388 2036 5396 2044
rect 5468 2036 5476 2044
rect 5532 2036 5540 2044
rect 6540 2036 6548 2044
rect 6668 2036 6676 2044
rect 7164 2036 7172 2044
rect 1411 2006 1419 2014
rect 1421 2006 1429 2014
rect 1431 2006 1439 2014
rect 1441 2006 1449 2014
rect 1451 2006 1459 2014
rect 1461 2006 1469 2014
rect 4419 2006 4427 2014
rect 4429 2006 4437 2014
rect 4439 2006 4447 2014
rect 4449 2006 4457 2014
rect 4459 2006 4467 2014
rect 4469 2006 4477 2014
rect 12 1976 20 1984
rect 188 1976 196 1984
rect 348 1976 356 1984
rect 556 1976 564 1984
rect 588 1976 596 1984
rect 652 1976 660 1984
rect 780 1976 788 1984
rect 940 1976 948 1984
rect 1324 1976 1332 1984
rect 1564 1976 1572 1984
rect 1596 1976 1604 1984
rect 1804 1976 1812 1984
rect 2188 1976 2196 1984
rect 2236 1976 2244 1984
rect 2668 1976 2676 1984
rect 2764 1976 2772 1984
rect 3356 1976 3364 1984
rect 3676 1976 3684 1984
rect 4060 1976 4068 1984
rect 4220 1976 4228 1984
rect 4252 1976 4260 1984
rect 4332 1976 4340 1984
rect 4508 1976 4516 1984
rect 4796 1976 4804 1984
rect 4860 1976 4868 1984
rect 4908 1976 4916 1984
rect 6124 1976 6132 1984
rect 6380 1976 6388 1984
rect 6540 1976 6548 1984
rect 6620 1976 6628 1984
rect 492 1956 500 1964
rect 4188 1956 4196 1964
rect 444 1936 452 1944
rect 508 1936 516 1944
rect 668 1936 676 1944
rect 940 1936 948 1944
rect 956 1936 964 1944
rect 1020 1936 1028 1944
rect 1116 1936 1124 1944
rect 1196 1936 1204 1944
rect 1308 1936 1316 1944
rect 1324 1936 1332 1944
rect 1372 1936 1380 1944
rect 1516 1936 1524 1944
rect 1548 1936 1556 1944
rect 1612 1936 1620 1944
rect 1676 1936 1684 1944
rect 1836 1936 1844 1944
rect 1900 1936 1908 1944
rect 1964 1936 1972 1944
rect 2076 1936 2084 1944
rect 2396 1936 2404 1944
rect 2460 1936 2468 1944
rect 2540 1936 2548 1944
rect 2812 1936 2820 1944
rect 3244 1936 3252 1944
rect 4172 1936 4180 1944
rect 4396 1936 4404 1944
rect 4652 1936 4660 1944
rect 4732 1936 4740 1944
rect 4780 1936 4788 1944
rect 5676 1936 5684 1944
rect 6476 1936 6484 1944
rect 204 1916 212 1924
rect 268 1916 276 1924
rect 396 1916 404 1924
rect 412 1916 420 1924
rect 476 1916 484 1924
rect 700 1916 708 1924
rect 924 1916 932 1924
rect 988 1916 996 1924
rect 1052 1916 1060 1924
rect 1164 1916 1172 1924
rect 1228 1916 1236 1924
rect 1340 1916 1348 1924
rect 1404 1916 1412 1924
rect 1484 1916 1492 1924
rect 1580 1916 1588 1924
rect 1644 1916 1652 1924
rect 1708 1916 1716 1924
rect 1868 1916 1876 1924
rect 1932 1916 1940 1924
rect 1996 1916 2004 1924
rect 2012 1916 2020 1924
rect 2108 1916 2116 1924
rect 2124 1916 2132 1924
rect 2284 1916 2292 1924
rect 2428 1916 2436 1924
rect 2476 1916 2484 1924
rect 2540 1916 2548 1924
rect 2604 1916 2612 1924
rect 2860 1916 2868 1924
rect 2892 1916 2900 1924
rect 2924 1916 2932 1924
rect 3052 1916 3060 1924
rect 3212 1916 3220 1924
rect 3276 1916 3284 1924
rect 3388 1916 3396 1924
rect 3500 1916 3508 1924
rect 3660 1916 3668 1924
rect 3852 1916 3860 1924
rect 3868 1916 3876 1924
rect 3932 1916 3940 1924
rect 3996 1916 4004 1924
rect 4092 1916 4100 1924
rect 4204 1916 4212 1924
rect 4284 1916 4292 1924
rect 4380 1916 4388 1924
rect 4428 1916 4436 1924
rect 4668 1916 4676 1924
rect 4764 1916 4772 1924
rect 5148 1916 5156 1924
rect 12 1896 20 1904
rect 108 1896 116 1904
rect 140 1896 148 1904
rect 172 1896 180 1904
rect 252 1896 260 1904
rect 284 1896 292 1904
rect 396 1896 404 1904
rect 428 1896 436 1904
rect 492 1896 500 1904
rect 572 1896 580 1904
rect 620 1896 628 1904
rect 684 1896 692 1904
rect 716 1896 724 1904
rect 876 1896 884 1904
rect 940 1896 948 1904
rect 1004 1896 1012 1904
rect 1068 1896 1076 1904
rect 1212 1896 1220 1904
rect 1260 1896 1268 1904
rect 1276 1896 1284 1904
rect 1324 1896 1332 1904
rect 1388 1896 1396 1904
rect 1564 1896 1572 1904
rect 1628 1896 1636 1904
rect 1692 1896 1700 1904
rect 1740 1896 1748 1904
rect 1788 1896 1796 1904
rect 1852 1896 1860 1904
rect 1916 1896 1924 1904
rect 1980 1896 1988 1904
rect 2012 1896 2020 1904
rect 2092 1896 2100 1904
rect 2124 1896 2132 1904
rect 2204 1896 2212 1904
rect 2268 1896 2276 1904
rect 2284 1896 2292 1904
rect 2316 1896 2324 1904
rect 2380 1896 2388 1904
rect 2492 1896 2500 1904
rect 2556 1896 2564 1904
rect 2732 1896 2740 1904
rect 172 1876 180 1884
rect 364 1876 372 1884
rect 636 1876 644 1884
rect 844 1880 852 1888
rect 44 1856 52 1864
rect 60 1856 68 1864
rect 108 1856 116 1864
rect 316 1856 324 1864
rect 332 1856 340 1864
rect 428 1856 436 1864
rect 540 1856 548 1864
rect 748 1856 756 1864
rect 860 1876 868 1884
rect 1052 1876 1060 1884
rect 1116 1876 1124 1884
rect 1132 1880 1140 1888
rect 1516 1876 1524 1884
rect 1692 1876 1700 1884
rect 1724 1876 1732 1884
rect 1916 1876 1924 1884
rect 2044 1876 2052 1884
rect 2156 1876 2164 1884
rect 2268 1876 2276 1884
rect 2460 1876 2468 1884
rect 2732 1876 2740 1884
rect 1212 1856 1220 1864
rect 1244 1856 1252 1864
rect 1788 1856 1796 1864
rect 1980 1856 1988 1864
rect 2172 1856 2180 1864
rect 2220 1856 2228 1864
rect 252 1836 260 1844
rect 364 1836 372 1844
rect 1852 1836 1860 1844
rect 2044 1836 2052 1844
rect 2076 1836 2084 1844
rect 2156 1836 2164 1844
rect 2412 1856 2420 1864
rect 2428 1856 2436 1864
rect 2604 1856 2612 1864
rect 2780 1896 2788 1904
rect 2860 1896 2868 1904
rect 2892 1896 2900 1904
rect 3020 1896 3028 1904
rect 3084 1896 3092 1904
rect 3180 1896 3188 1904
rect 3244 1896 3252 1904
rect 3308 1896 3316 1904
rect 3420 1896 3428 1904
rect 3452 1896 3460 1904
rect 3580 1896 3588 1904
rect 2908 1876 2916 1884
rect 3036 1876 3044 1884
rect 3100 1876 3108 1884
rect 3196 1876 3204 1884
rect 3260 1876 3268 1884
rect 3324 1876 3332 1884
rect 3404 1876 3412 1884
rect 3468 1876 3476 1884
rect 3548 1876 3556 1884
rect 3612 1876 3620 1884
rect 3692 1876 3700 1884
rect 3740 1876 3748 1884
rect 3820 1896 3828 1904
rect 3916 1896 3924 1904
rect 3948 1896 3956 1904
rect 3996 1896 4004 1904
rect 4012 1896 4020 1904
rect 4028 1896 4036 1904
rect 4076 1896 4084 1904
rect 4124 1896 4132 1904
rect 4188 1896 4196 1904
rect 4364 1896 4372 1904
rect 4412 1896 4420 1904
rect 4748 1896 4756 1904
rect 4796 1896 4804 1904
rect 5004 1896 5012 1904
rect 5052 1896 5060 1904
rect 5148 1896 5156 1904
rect 5196 1916 5204 1924
rect 5708 1916 5716 1924
rect 5740 1916 5748 1924
rect 6236 1916 6244 1924
rect 6444 1916 6452 1924
rect 6604 1916 6612 1924
rect 6860 1916 6868 1924
rect 6924 1916 6932 1924
rect 6956 1916 6964 1924
rect 5276 1896 5284 1904
rect 5340 1896 5348 1904
rect 5452 1896 5460 1904
rect 5580 1896 5588 1904
rect 5644 1896 5652 1904
rect 5676 1896 5684 1904
rect 5756 1896 5764 1904
rect 5772 1896 5780 1904
rect 5788 1896 5796 1904
rect 5852 1896 5860 1904
rect 5884 1896 5892 1904
rect 5916 1896 5924 1904
rect 6012 1896 6020 1904
rect 6028 1896 6036 1904
rect 6092 1896 6100 1904
rect 6140 1896 6148 1904
rect 6188 1896 6196 1904
rect 6284 1896 6292 1904
rect 6316 1896 6324 1904
rect 6428 1896 6436 1904
rect 6572 1896 6580 1904
rect 6684 1896 6692 1904
rect 6732 1896 6740 1904
rect 6844 1896 6852 1904
rect 6908 1896 6916 1904
rect 6956 1896 6964 1904
rect 7100 1896 7108 1904
rect 7244 1896 7252 1904
rect 7308 1894 7316 1902
rect 3772 1876 3780 1884
rect 3804 1876 3812 1884
rect 3836 1876 3844 1884
rect 3868 1876 3876 1884
rect 3980 1876 3988 1884
rect 4044 1876 4052 1884
rect 4140 1876 4148 1884
rect 4316 1876 4324 1884
rect 2812 1856 2820 1864
rect 2844 1856 2852 1864
rect 3132 1856 3140 1864
rect 3644 1856 3652 1864
rect 3708 1856 3716 1864
rect 3772 1856 3780 1864
rect 4076 1856 4084 1864
rect 4236 1856 4244 1864
rect 4268 1856 4276 1864
rect 4300 1856 4308 1864
rect 4620 1876 4628 1884
rect 4700 1876 4708 1884
rect 4844 1876 4852 1884
rect 4892 1876 4900 1884
rect 4956 1876 4964 1884
rect 5132 1876 5140 1884
rect 5228 1876 5236 1884
rect 5324 1876 5332 1884
rect 5420 1876 5428 1884
rect 5580 1876 5588 1884
rect 5628 1876 5636 1884
rect 5644 1876 5652 1884
rect 5852 1876 5860 1884
rect 5900 1876 5908 1884
rect 5932 1876 5940 1884
rect 6412 1876 6420 1884
rect 6476 1876 6484 1884
rect 6492 1876 6500 1884
rect 6508 1880 6516 1888
rect 6556 1876 6564 1884
rect 6652 1876 6660 1884
rect 6892 1876 6900 1884
rect 6972 1876 6980 1884
rect 7116 1876 7124 1884
rect 4540 1856 4548 1864
rect 4556 1856 4564 1864
rect 4604 1856 4612 1864
rect 5244 1856 5252 1864
rect 5308 1856 5316 1864
rect 5548 1856 5556 1864
rect 5724 1856 5732 1864
rect 6044 1856 6052 1864
rect 6108 1856 6116 1864
rect 6156 1856 6164 1864
rect 6204 1856 6212 1864
rect 6220 1856 6228 1864
rect 6284 1856 6292 1864
rect 6348 1856 6356 1864
rect 6364 1856 6372 1864
rect 6396 1856 6404 1864
rect 6812 1856 6820 1864
rect 2524 1836 2532 1844
rect 2620 1836 2628 1844
rect 2988 1836 2996 1844
rect 3052 1836 3060 1844
rect 3148 1836 3156 1844
rect 3276 1836 3284 1844
rect 3724 1836 3732 1844
rect 3788 1836 3796 1844
rect 5116 1836 5124 1844
rect 5532 1836 5540 1844
rect 5804 1836 5812 1844
rect 6172 1836 6180 1844
rect 6300 1836 6308 1844
rect 6460 1836 6468 1844
rect 6604 1836 6612 1844
rect 6988 1836 6996 1844
rect 7180 1836 7188 1844
rect 60 1816 68 1824
rect 2915 1806 2923 1814
rect 2925 1806 2933 1814
rect 2935 1806 2943 1814
rect 2945 1806 2953 1814
rect 2955 1806 2963 1814
rect 2965 1806 2973 1814
rect 5923 1806 5931 1814
rect 5933 1806 5941 1814
rect 5943 1806 5951 1814
rect 5953 1806 5961 1814
rect 5963 1806 5971 1814
rect 5973 1806 5981 1814
rect 12 1796 20 1804
rect 124 1796 132 1804
rect 380 1796 388 1804
rect 508 1796 516 1804
rect 1244 1796 1252 1804
rect 2044 1796 2052 1804
rect 2156 1796 2164 1804
rect 2268 1796 2276 1804
rect 2652 1796 2660 1804
rect 60 1776 68 1784
rect 396 1776 404 1784
rect 588 1776 596 1784
rect 700 1776 708 1784
rect 716 1776 724 1784
rect 972 1776 980 1784
rect 1068 1776 1076 1784
rect 12 1756 20 1764
rect 124 1756 132 1764
rect 236 1756 244 1764
rect 268 1756 276 1764
rect 380 1756 388 1764
rect 412 1756 420 1764
rect 476 1756 484 1764
rect 508 1756 516 1764
rect 540 1756 548 1764
rect 572 1756 580 1764
rect 876 1756 884 1764
rect 1052 1756 1060 1764
rect 1292 1776 1300 1784
rect 1372 1776 1380 1784
rect 1148 1756 1156 1764
rect 108 1736 116 1744
rect 188 1736 196 1744
rect 236 1736 244 1744
rect 268 1736 276 1744
rect 428 1736 436 1744
rect 636 1736 644 1744
rect 764 1736 772 1744
rect 780 1736 788 1744
rect 860 1736 868 1744
rect 940 1736 948 1744
rect 1036 1736 1044 1744
rect 1244 1756 1252 1764
rect 1356 1756 1364 1764
rect 1516 1776 1524 1784
rect 1836 1776 1844 1784
rect 2108 1776 2116 1784
rect 2220 1776 2228 1784
rect 2284 1776 2292 1784
rect 1580 1756 1588 1764
rect 1244 1736 1252 1744
rect 1340 1736 1348 1744
rect 1564 1736 1572 1744
rect 1628 1756 1636 1764
rect 1740 1756 1748 1764
rect 1676 1736 1684 1744
rect 1788 1756 1796 1764
rect 1996 1756 2004 1764
rect 2044 1756 2052 1764
rect 2156 1756 2164 1764
rect 2268 1756 2276 1764
rect 2332 1756 2340 1764
rect 2476 1776 2484 1784
rect 2524 1776 2532 1784
rect 2668 1776 2676 1784
rect 2828 1776 2836 1784
rect 2876 1776 2884 1784
rect 3340 1776 3348 1784
rect 3388 1776 3396 1784
rect 3436 1776 3444 1784
rect 3708 1776 3716 1784
rect 3772 1776 3780 1784
rect 3980 1776 3988 1784
rect 4012 1776 4020 1784
rect 4044 1776 4052 1784
rect 4092 1776 4100 1784
rect 4220 1776 4228 1784
rect 4332 1776 4340 1784
rect 4492 1776 4500 1784
rect 4668 1776 4676 1784
rect 4844 1776 4852 1784
rect 5020 1776 5028 1784
rect 5228 1776 5236 1784
rect 6268 1776 6276 1784
rect 6652 1776 6660 1784
rect 6764 1776 6772 1784
rect 2492 1756 2500 1764
rect 2508 1756 2516 1764
rect 2652 1756 2660 1764
rect 1884 1736 1892 1744
rect 1948 1736 1956 1744
rect 2044 1736 2052 1744
rect 2156 1736 2164 1744
rect 2316 1736 2324 1744
rect 2332 1736 2340 1744
rect 2540 1736 2548 1744
rect 2716 1736 2724 1744
rect 2764 1756 2772 1764
rect 3500 1756 3508 1764
rect 4028 1756 4036 1764
rect 4060 1756 4068 1764
rect 4124 1756 4132 1764
rect 4140 1756 4148 1764
rect 4188 1756 4196 1764
rect 4252 1756 4260 1764
rect 4284 1756 4292 1764
rect 4316 1756 4324 1764
rect 4556 1756 4564 1764
rect 4572 1756 4580 1764
rect 4620 1756 4628 1764
rect 4828 1756 4836 1764
rect 4892 1756 4900 1764
rect 5420 1756 5428 1764
rect 5532 1756 5540 1764
rect 5724 1756 5732 1764
rect 5740 1756 5748 1764
rect 6204 1756 6212 1764
rect 6316 1756 6324 1764
rect 6412 1756 6420 1764
rect 6540 1756 6548 1764
rect 6636 1756 6644 1764
rect 6860 1756 6868 1764
rect 7036 1756 7044 1764
rect 2780 1736 2788 1744
rect 2844 1736 2852 1744
rect 2940 1736 2948 1744
rect 3228 1736 3236 1744
rect 3260 1736 3268 1744
rect 3356 1736 3364 1744
rect 3756 1736 3764 1744
rect 3820 1736 3828 1744
rect 3836 1736 3844 1744
rect 3932 1736 3940 1744
rect 3964 1736 3972 1744
rect 4076 1736 4084 1744
rect 4204 1736 4212 1744
rect 4540 1736 4548 1744
rect 4716 1736 4724 1744
rect 60 1716 68 1724
rect 92 1716 100 1724
rect 172 1716 180 1724
rect 204 1716 212 1724
rect 284 1716 292 1724
rect 300 1716 308 1724
rect 332 1716 340 1724
rect 428 1716 436 1724
rect 476 1716 484 1724
rect 540 1716 548 1724
rect 620 1716 628 1724
rect 668 1716 676 1724
rect 748 1716 756 1724
rect 812 1716 820 1724
rect 924 1716 932 1724
rect 1084 1716 1092 1724
rect 1148 1716 1156 1724
rect 1180 1716 1188 1724
rect 1292 1716 1300 1724
rect 1324 1716 1332 1724
rect 1388 1716 1396 1724
rect 1516 1716 1524 1724
rect 1548 1716 1556 1724
rect 1580 1716 1588 1724
rect 1660 1716 1668 1724
rect 1692 1716 1700 1724
rect 1820 1716 1828 1724
rect 1868 1716 1876 1724
rect 1948 1716 1956 1724
rect 1964 1716 1972 1724
rect 1996 1716 2004 1724
rect 2060 1716 2068 1724
rect 2108 1716 2116 1724
rect 2188 1716 2196 1724
rect 2220 1716 2228 1724
rect 2364 1716 2372 1724
rect 2396 1716 2404 1724
rect 2460 1716 2468 1724
rect 2540 1716 2548 1724
rect 2572 1716 2580 1724
rect 2604 1716 2612 1724
rect 2700 1716 2708 1724
rect 2764 1716 2772 1724
rect 2796 1716 2804 1724
rect 3196 1718 3204 1726
rect 3276 1716 3284 1724
rect 3372 1716 3380 1724
rect 3420 1716 3428 1724
rect 3468 1716 3476 1724
rect 3596 1716 3604 1724
rect 3644 1718 3652 1726
rect 3740 1716 3748 1724
rect 3804 1716 3812 1724
rect 3916 1716 3924 1724
rect 3948 1716 3956 1724
rect 300 1696 308 1704
rect 828 1696 836 1704
rect 1436 1696 1444 1704
rect 1484 1696 1492 1704
rect 2396 1696 2404 1704
rect 2572 1696 2580 1704
rect 3308 1696 3316 1704
rect 3708 1696 3716 1704
rect 3772 1696 3780 1704
rect 3884 1696 3892 1704
rect 3996 1696 4004 1704
rect 4108 1696 4116 1704
rect 4476 1716 4484 1724
rect 4524 1716 4532 1724
rect 4620 1716 4628 1724
rect 4780 1736 4788 1744
rect 4828 1736 4836 1744
rect 4908 1736 4916 1744
rect 4940 1736 4948 1744
rect 4988 1736 4996 1744
rect 5036 1736 5044 1744
rect 5068 1736 5076 1744
rect 5244 1736 5252 1744
rect 5276 1736 5284 1744
rect 5308 1736 5316 1744
rect 5372 1736 5380 1744
rect 5580 1736 5588 1744
rect 5644 1736 5652 1744
rect 5660 1736 5668 1744
rect 5772 1736 5780 1744
rect 5836 1736 5844 1744
rect 5852 1736 5860 1744
rect 5884 1736 5892 1744
rect 6220 1736 6228 1744
rect 6300 1736 6308 1744
rect 6364 1736 6372 1744
rect 6428 1736 6436 1744
rect 6492 1736 6500 1744
rect 6556 1736 6564 1744
rect 6620 1736 6628 1744
rect 6684 1736 6692 1744
rect 6732 1736 6740 1744
rect 6748 1736 6756 1744
rect 6812 1736 6820 1744
rect 6860 1736 6868 1744
rect 6908 1736 6916 1744
rect 7004 1736 7012 1744
rect 7036 1736 7044 1744
rect 7052 1736 7060 1744
rect 7148 1736 7156 1744
rect 4780 1716 4788 1724
rect 4684 1696 4692 1704
rect 4764 1696 4772 1704
rect 5132 1716 5140 1724
rect 5260 1716 5268 1724
rect 5324 1716 5332 1724
rect 5340 1716 5348 1724
rect 5372 1716 5380 1724
rect 5388 1716 5396 1724
rect 5452 1716 5460 1724
rect 5500 1716 5508 1724
rect 5516 1716 5524 1724
rect 5564 1716 5572 1724
rect 5596 1716 5604 1724
rect 5644 1716 5652 1724
rect 5676 1716 5684 1724
rect 5756 1716 5764 1724
rect 5788 1716 5796 1724
rect 5820 1716 5828 1724
rect 5868 1716 5876 1724
rect 5996 1716 6004 1724
rect 6044 1716 6052 1724
rect 6060 1716 6068 1724
rect 6092 1716 6100 1724
rect 6140 1716 6148 1724
rect 6156 1716 6164 1724
rect 6172 1716 6180 1724
rect 6300 1716 6308 1724
rect 6348 1716 6356 1724
rect 6380 1716 6388 1724
rect 6444 1716 6452 1724
rect 6492 1716 6500 1724
rect 6508 1716 6516 1724
rect 6572 1716 6580 1724
rect 6604 1716 6612 1724
rect 6668 1716 6676 1724
rect 6700 1716 6708 1724
rect 4940 1696 4948 1704
rect 5292 1696 5300 1704
rect 5676 1696 5684 1704
rect 5708 1696 5716 1704
rect 5900 1696 5908 1704
rect 6252 1696 6260 1704
rect 6268 1696 6276 1704
rect 6412 1696 6420 1704
rect 6764 1716 6772 1724
rect 6812 1716 6820 1724
rect 6828 1716 6836 1724
rect 6892 1716 6900 1724
rect 6972 1716 6980 1724
rect 6988 1716 6996 1724
rect 6924 1696 6932 1704
rect 7084 1696 7092 1704
rect 7132 1716 7140 1724
rect 7244 1716 7252 1724
rect 7276 1716 7284 1724
rect 7132 1696 7140 1704
rect 1884 1676 1892 1684
rect 3100 1676 3108 1684
rect 3500 1676 3508 1684
rect 3516 1676 3524 1684
rect 5388 1676 5396 1684
rect 6508 1676 6516 1684
rect 6828 1676 6836 1684
rect 7164 1676 7172 1684
rect 4380 1656 4388 1664
rect 5820 1656 5828 1664
rect 2956 1636 2964 1644
rect 3068 1636 3076 1644
rect 4572 1636 4580 1644
rect 4972 1636 4980 1644
rect 5468 1636 5476 1644
rect 5564 1636 5572 1644
rect 5596 1636 5604 1644
rect 6012 1636 6020 1644
rect 6108 1636 6116 1644
rect 6236 1636 6244 1644
rect 6284 1636 6292 1644
rect 6444 1636 6452 1644
rect 6572 1636 6580 1644
rect 6940 1636 6948 1644
rect 1411 1606 1419 1614
rect 1421 1606 1429 1614
rect 1431 1606 1439 1614
rect 1441 1606 1449 1614
rect 1451 1606 1459 1614
rect 1461 1606 1469 1614
rect 4419 1606 4427 1614
rect 4429 1606 4437 1614
rect 4439 1606 4447 1614
rect 4449 1606 4457 1614
rect 4459 1606 4467 1614
rect 4469 1606 4477 1614
rect 28 1576 36 1584
rect 60 1576 68 1584
rect 124 1576 132 1584
rect 156 1576 164 1584
rect 220 1576 228 1584
rect 284 1576 292 1584
rect 700 1576 708 1584
rect 764 1576 772 1584
rect 1084 1576 1092 1584
rect 1260 1576 1268 1584
rect 1356 1576 1364 1584
rect 1484 1576 1492 1584
rect 1676 1576 1684 1584
rect 1916 1576 1924 1584
rect 2012 1576 2020 1584
rect 2124 1576 2132 1584
rect 2220 1576 2228 1584
rect 2316 1576 2324 1584
rect 2348 1576 2356 1584
rect 2556 1576 2564 1584
rect 2620 1576 2628 1584
rect 2828 1576 2836 1584
rect 3644 1576 3652 1584
rect 3964 1576 3972 1584
rect 4012 1576 4020 1584
rect 4124 1576 4132 1584
rect 4316 1576 4324 1584
rect 4380 1576 4388 1584
rect 4556 1576 4564 1584
rect 4636 1576 4644 1584
rect 4716 1576 4724 1584
rect 4748 1576 4756 1584
rect 4812 1576 4820 1584
rect 4876 1576 4884 1584
rect 5884 1576 5892 1584
rect 6204 1576 6212 1584
rect 6524 1576 6532 1584
rect 6604 1576 6612 1584
rect 6700 1576 6708 1584
rect 7180 1576 7188 1584
rect 7276 1576 7284 1584
rect 7356 1576 7364 1584
rect 2940 1556 2948 1564
rect 3852 1556 3860 1564
rect 684 1536 692 1544
rect 780 1536 788 1544
rect 1068 1536 1076 1544
rect 1148 1536 1156 1544
rect 1228 1536 1236 1544
rect 3836 1536 3844 1544
rect 3996 1536 4004 1544
rect 4044 1536 4052 1544
rect 4108 1536 4116 1544
rect 4268 1536 4276 1544
rect 4332 1536 4340 1544
rect 4396 1536 4404 1544
rect 4620 1536 4628 1544
rect 4652 1536 4660 1544
rect 4700 1536 4708 1544
rect 4764 1536 4772 1544
rect 4828 1536 4836 1544
rect 6268 1536 6276 1544
rect 6764 1536 6772 1544
rect 636 1516 644 1524
rect 684 1516 692 1524
rect 748 1516 756 1524
rect 844 1516 852 1524
rect 204 1496 212 1504
rect 284 1496 292 1504
rect 316 1496 324 1504
rect 348 1496 356 1504
rect 364 1496 372 1504
rect 76 1476 84 1484
rect 92 1480 100 1488
rect 300 1476 308 1484
rect 396 1476 404 1484
rect 540 1496 548 1504
rect 700 1496 708 1504
rect 764 1496 772 1504
rect 1100 1516 1108 1524
rect 1596 1516 1604 1524
rect 1836 1516 1844 1524
rect 2812 1516 2820 1524
rect 3244 1516 3252 1524
rect 3324 1516 3332 1524
rect 892 1496 900 1504
rect 924 1496 932 1504
rect 1036 1496 1044 1504
rect 1084 1496 1092 1504
rect 1388 1496 1396 1504
rect 1516 1496 1524 1504
rect 1564 1496 1572 1504
rect 1724 1496 1732 1504
rect 1788 1496 1796 1504
rect 1804 1496 1812 1504
rect 1868 1496 1876 1504
rect 1948 1496 1956 1504
rect 2044 1496 2052 1504
rect 2076 1496 2084 1504
rect 2380 1496 2388 1504
rect 2428 1496 2436 1504
rect 2460 1496 2468 1504
rect 2524 1496 2532 1504
rect 2556 1496 2564 1504
rect 2588 1496 2596 1504
rect 2652 1496 2660 1504
rect 2700 1496 2708 1504
rect 2860 1496 2868 1504
rect 3036 1496 3044 1504
rect 3196 1496 3204 1504
rect 3212 1496 3220 1504
rect 3308 1496 3316 1504
rect 3356 1496 3364 1504
rect 3436 1496 3444 1504
rect 3484 1496 3492 1504
rect 3500 1496 3508 1504
rect 3564 1516 3572 1524
rect 3660 1516 3668 1524
rect 3708 1516 3716 1524
rect 3804 1516 3812 1524
rect 3868 1516 3876 1524
rect 3884 1516 3892 1524
rect 4028 1516 4036 1524
rect 4140 1516 4148 1524
rect 4156 1516 4164 1524
rect 4300 1516 4308 1524
rect 4364 1516 4372 1524
rect 4428 1516 4436 1524
rect 4588 1516 4596 1524
rect 4620 1516 4628 1524
rect 4732 1516 4740 1524
rect 4796 1516 4804 1524
rect 4860 1516 4868 1524
rect 6364 1516 6372 1524
rect 6988 1516 6996 1524
rect 3612 1496 3620 1504
rect 3740 1496 3748 1504
rect 3852 1496 3860 1504
rect 3932 1496 3940 1504
rect 4012 1496 4020 1504
rect 4124 1496 4132 1504
rect 492 1476 500 1484
rect 556 1476 564 1484
rect 572 1476 580 1484
rect 668 1476 676 1484
rect 812 1476 820 1484
rect 908 1476 916 1484
rect 972 1476 980 1484
rect 1212 1476 1220 1484
rect 1324 1476 1332 1484
rect 1500 1476 1508 1484
rect 1564 1476 1572 1484
rect 1612 1476 1620 1484
rect 1740 1476 1748 1484
rect 1900 1476 1908 1484
rect 1932 1476 1940 1484
rect 2156 1476 2164 1484
rect 2252 1476 2260 1484
rect 2364 1476 2372 1484
rect 2476 1476 2484 1484
rect 2492 1480 2500 1488
rect 2540 1476 2548 1484
rect 2604 1476 2612 1484
rect 2668 1476 2676 1484
rect 2748 1476 2756 1484
rect 3100 1476 3108 1484
rect 3164 1476 3172 1484
rect 3196 1476 3204 1484
rect 3292 1476 3300 1484
rect 3340 1476 3348 1484
rect 3372 1476 3380 1484
rect 3420 1476 3428 1484
rect 3500 1476 3508 1484
rect 3532 1476 3540 1484
rect 3596 1476 3604 1484
rect 3676 1476 3684 1484
rect 3692 1476 3700 1484
rect 3756 1476 3764 1484
rect 3788 1476 3796 1484
rect 3916 1476 3924 1484
rect 4076 1476 4084 1484
rect 4188 1476 4196 1484
rect 4284 1496 4292 1504
rect 4348 1496 4356 1504
rect 4412 1496 4420 1504
rect 4588 1496 4596 1504
rect 4636 1496 4644 1504
rect 4716 1496 4724 1504
rect 4780 1496 4788 1504
rect 4844 1496 4852 1504
rect 4988 1496 4996 1504
rect 5100 1496 5108 1504
rect 5212 1496 5220 1504
rect 5228 1496 5236 1504
rect 5276 1496 5284 1504
rect 5292 1496 5300 1504
rect 5308 1496 5316 1504
rect 5372 1496 5380 1504
rect 5420 1496 5428 1504
rect 5468 1496 5476 1504
rect 5516 1496 5524 1504
rect 5644 1496 5652 1504
rect 5692 1496 5700 1504
rect 5804 1496 5812 1504
rect 5868 1496 5876 1504
rect 5916 1496 5924 1504
rect 5996 1496 6004 1504
rect 6044 1496 6052 1504
rect 6092 1496 6100 1504
rect 6140 1496 6148 1504
rect 6204 1496 6212 1504
rect 6252 1496 6260 1504
rect 6268 1496 6276 1504
rect 6332 1496 6340 1504
rect 6396 1496 6404 1504
rect 6444 1496 6452 1504
rect 6460 1496 6468 1504
rect 6476 1496 6484 1504
rect 6492 1496 6500 1504
rect 6556 1496 6564 1504
rect 6588 1496 6596 1504
rect 6636 1496 6644 1504
rect 6652 1496 6660 1504
rect 6684 1496 6692 1504
rect 6732 1496 6740 1504
rect 6748 1496 6756 1504
rect 7340 1516 7348 1524
rect 6892 1494 6900 1502
rect 7036 1496 7044 1504
rect 7068 1496 7076 1504
rect 7132 1496 7140 1504
rect 7164 1496 7172 1504
rect 7180 1496 7188 1504
rect 7228 1496 7236 1504
rect 7292 1496 7300 1504
rect 4508 1476 4516 1484
rect 4956 1476 4964 1484
rect 5116 1476 5124 1484
rect 12 1456 20 1464
rect 44 1456 52 1464
rect 140 1456 148 1464
rect 172 1456 180 1464
rect 188 1456 196 1464
rect 236 1456 244 1464
rect 252 1456 260 1464
rect 444 1456 452 1464
rect 460 1456 468 1464
rect 844 1456 852 1464
rect 924 1456 932 1464
rect 956 1456 964 1464
rect 972 1456 980 1464
rect 1036 1456 1044 1464
rect 1228 1456 1236 1464
rect 1340 1456 1348 1464
rect 1372 1456 1380 1464
rect 1788 1456 1796 1464
rect 1820 1456 1828 1464
rect 1900 1456 1908 1464
rect 2076 1456 2084 1464
rect 2140 1456 2148 1464
rect 2236 1456 2244 1464
rect 2300 1456 2308 1464
rect 2332 1456 2340 1464
rect 2428 1456 2436 1464
rect 2444 1456 2452 1464
rect 2668 1456 2676 1464
rect 2764 1456 2772 1464
rect 3132 1456 3140 1464
rect 3388 1456 3396 1464
rect 4044 1456 4052 1464
rect 4236 1456 4244 1464
rect 4524 1456 4532 1464
rect 4892 1456 4900 1464
rect 5324 1476 5332 1484
rect 5516 1476 5524 1484
rect 5532 1476 5540 1484
rect 5564 1476 5572 1484
rect 5852 1476 5860 1484
rect 6124 1476 6132 1484
rect 6188 1476 6196 1484
rect 6252 1476 6260 1484
rect 6316 1476 6324 1484
rect 6348 1476 6356 1484
rect 6380 1476 6388 1484
rect 6924 1476 6932 1484
rect 6956 1476 6964 1484
rect 7052 1476 7060 1484
rect 7084 1476 7092 1484
rect 5164 1456 5172 1464
rect 5404 1456 5412 1464
rect 5500 1456 5508 1464
rect 5564 1456 5572 1464
rect 5772 1456 5780 1464
rect 6300 1456 6308 1464
rect 7244 1476 7252 1484
rect 7372 1476 7380 1484
rect 7132 1456 7140 1464
rect 7212 1456 7220 1464
rect 7324 1456 7332 1464
rect 428 1436 436 1444
rect 508 1436 516 1444
rect 860 1436 868 1444
rect 1548 1436 1556 1444
rect 1756 1436 1764 1444
rect 2284 1436 2292 1444
rect 2716 1436 2724 1444
rect 2796 1436 2804 1444
rect 3148 1436 3156 1444
rect 3276 1436 3284 1444
rect 3404 1436 3412 1444
rect 3708 1436 3716 1444
rect 3900 1436 3908 1444
rect 5084 1436 5092 1444
rect 5132 1436 5140 1444
rect 5244 1436 5252 1444
rect 5340 1436 5348 1444
rect 5452 1436 5460 1444
rect 5580 1436 5588 1444
rect 5836 1436 5844 1444
rect 5884 1436 5892 1444
rect 6028 1436 6036 1444
rect 6076 1436 6084 1444
rect 6172 1436 6180 1444
rect 7004 1436 7012 1444
rect 2915 1406 2923 1414
rect 2925 1406 2933 1414
rect 2935 1406 2943 1414
rect 2945 1406 2953 1414
rect 2955 1406 2963 1414
rect 2965 1406 2973 1414
rect 5923 1406 5931 1414
rect 5933 1406 5941 1414
rect 5943 1406 5951 1414
rect 5953 1406 5961 1414
rect 5963 1406 5971 1414
rect 5973 1406 5981 1414
rect 12 1376 20 1384
rect 412 1376 420 1384
rect 652 1376 660 1384
rect 716 1376 724 1384
rect 748 1376 756 1384
rect 876 1376 884 1384
rect 940 1376 948 1384
rect 1004 1376 1012 1384
rect 1084 1376 1092 1384
rect 1212 1376 1220 1384
rect 1516 1376 1524 1384
rect 1564 1376 1572 1384
rect 1708 1376 1716 1384
rect 2012 1376 2020 1384
rect 2204 1376 2212 1384
rect 2300 1376 2308 1384
rect 2364 1376 2372 1384
rect 2412 1376 2420 1384
rect 2524 1376 2532 1384
rect 2604 1376 2612 1384
rect 2716 1376 2724 1384
rect 3004 1376 3012 1384
rect 3420 1376 3428 1384
rect 3772 1376 3780 1384
rect 3820 1376 3828 1384
rect 3948 1376 3956 1384
rect 4012 1376 4020 1384
rect 4156 1376 4164 1384
rect 4444 1376 4452 1384
rect 4812 1376 4820 1384
rect 5404 1376 5412 1384
rect 5708 1376 5716 1384
rect 6636 1376 6644 1384
rect 6732 1376 6740 1384
rect 7116 1376 7124 1384
rect 60 1356 68 1364
rect 140 1356 148 1364
rect 204 1356 212 1364
rect 268 1356 276 1364
rect 300 1356 308 1364
rect 316 1356 324 1364
rect 492 1356 500 1364
rect 508 1356 516 1364
rect 732 1356 740 1364
rect 1068 1356 1076 1364
rect 1180 1356 1188 1364
rect 1260 1356 1268 1364
rect 1324 1356 1332 1364
rect 1340 1356 1348 1364
rect 1548 1356 1556 1364
rect 1580 1356 1588 1364
rect 1836 1356 1844 1364
rect 1868 1356 1876 1364
rect 1884 1356 1892 1364
rect 1932 1356 1940 1364
rect 2028 1356 2036 1364
rect 2044 1356 2052 1364
rect 2156 1356 2164 1364
rect 2348 1356 2356 1364
rect 2620 1356 2628 1364
rect 3148 1356 3156 1364
rect 3628 1356 3636 1364
rect 3708 1356 3716 1364
rect 3740 1356 3748 1364
rect 3788 1356 3796 1364
rect 4028 1356 4036 1364
rect 4108 1356 4116 1364
rect 4172 1356 4180 1364
rect 4252 1356 4260 1364
rect 4684 1356 4692 1364
rect 5276 1356 5284 1364
rect 6412 1356 6420 1364
rect 6460 1356 6468 1364
rect 76 1336 84 1344
rect 332 1336 340 1344
rect 364 1336 372 1344
rect 460 1336 468 1344
rect 540 1336 548 1344
rect 636 1336 644 1344
rect 700 1336 708 1344
rect 844 1336 852 1344
rect 892 1336 900 1344
rect 1052 1336 1060 1344
rect 1100 1336 1108 1344
rect 1132 1336 1140 1344
rect 1212 1336 1220 1344
rect 1500 1336 1508 1344
rect 1532 1336 1540 1344
rect 1596 1336 1604 1344
rect 1660 1336 1668 1344
rect 1820 1336 1828 1344
rect 92 1316 100 1324
rect 124 1316 132 1324
rect 172 1316 180 1324
rect 220 1316 228 1324
rect 236 1316 244 1324
rect 284 1316 292 1324
rect 348 1316 356 1324
rect 492 1316 500 1324
rect 556 1316 564 1324
rect 604 1316 612 1324
rect 780 1316 788 1324
rect 796 1316 804 1324
rect 908 1316 916 1324
rect 1116 1316 1124 1324
rect 1180 1316 1188 1324
rect 1292 1316 1300 1324
rect 1308 1316 1316 1324
rect 1372 1316 1380 1324
rect 1548 1316 1556 1324
rect 1612 1316 1620 1324
rect 1804 1316 1812 1324
rect 1836 1316 1844 1324
rect 1996 1336 2004 1344
rect 2028 1336 2036 1344
rect 2124 1332 2132 1340
rect 2284 1336 2292 1344
rect 2332 1336 2340 1344
rect 1980 1316 1988 1324
rect 2076 1316 2084 1324
rect 2188 1316 2196 1324
rect 2396 1316 2404 1324
rect 2444 1316 2452 1324
rect 2556 1336 2564 1344
rect 2572 1336 2580 1344
rect 2604 1336 2612 1344
rect 2700 1336 2708 1344
rect 2732 1336 2740 1344
rect 2764 1336 2772 1344
rect 2860 1336 2868 1344
rect 2892 1336 2900 1344
rect 3212 1336 3220 1344
rect 3308 1336 3316 1344
rect 3324 1336 3332 1344
rect 3580 1336 3588 1344
rect 3868 1336 3876 1344
rect 3884 1332 3892 1340
rect 4188 1336 4196 1344
rect 4364 1336 4372 1344
rect 4828 1336 4836 1344
rect 4924 1336 4932 1344
rect 5900 1336 5908 1344
rect 6028 1336 6036 1344
rect 6060 1336 6068 1344
rect 6092 1336 6100 1344
rect 6220 1336 6228 1344
rect 6332 1336 6340 1344
rect 6364 1336 6372 1344
rect 6412 1336 6420 1344
rect 6476 1336 6484 1344
rect 6588 1336 6596 1344
rect 6796 1336 6804 1344
rect 6908 1336 6916 1344
rect 7052 1336 7060 1344
rect 7212 1336 7220 1344
rect 7340 1336 7348 1344
rect 2492 1316 2500 1324
rect 2748 1316 2756 1324
rect 2764 1316 2772 1324
rect 2876 1316 2884 1324
rect 2908 1316 2916 1324
rect 3148 1318 3156 1326
rect 3228 1316 3236 1324
rect 3324 1316 3332 1324
rect 3372 1316 3380 1324
rect 3388 1316 3396 1324
rect 3468 1316 3476 1324
rect 3516 1316 3524 1324
rect 3532 1316 3540 1324
rect 3596 1316 3604 1324
rect 3676 1316 3684 1324
rect 3836 1316 3844 1324
rect 3948 1316 3956 1324
rect 3996 1316 4004 1324
rect 4076 1316 4084 1324
rect 4508 1316 4516 1324
rect 4572 1318 4580 1326
rect 4700 1316 4708 1324
rect 620 1296 628 1304
rect 668 1296 676 1304
rect 892 1296 900 1304
rect 1212 1296 1220 1304
rect 1372 1296 1380 1304
rect 1404 1296 1412 1304
rect 1644 1296 1652 1304
rect 1772 1296 1780 1304
rect 1884 1296 1892 1304
rect 2172 1296 2180 1304
rect 2204 1296 2212 1304
rect 2252 1296 2260 1304
rect 2604 1296 2612 1304
rect 2812 1296 2820 1304
rect 2940 1296 2948 1304
rect 3260 1296 3268 1304
rect 3628 1296 3636 1304
rect 3852 1296 3860 1304
rect 3932 1296 3940 1304
rect 4044 1296 4052 1304
rect 4092 1296 4100 1304
rect 4860 1296 4868 1304
rect 4908 1316 4916 1324
rect 4988 1318 4996 1326
rect 5052 1316 5060 1324
rect 5164 1316 5172 1324
rect 5212 1316 5220 1324
rect 5324 1316 5332 1324
rect 5420 1316 5428 1324
rect 5436 1316 5444 1324
rect 5500 1316 5508 1324
rect 5516 1316 5524 1324
rect 5532 1316 5540 1324
rect 5580 1316 5588 1324
rect 5628 1316 5636 1324
rect 5676 1316 5684 1324
rect 5692 1316 5700 1324
rect 5772 1316 5780 1324
rect 5836 1318 5844 1326
rect 5916 1316 5924 1324
rect 6044 1316 6052 1324
rect 6108 1316 6116 1324
rect 6172 1316 6180 1324
rect 6204 1316 6212 1324
rect 6236 1316 6244 1324
rect 6316 1316 6324 1324
rect 6348 1316 6356 1324
rect 6380 1316 6388 1324
rect 6428 1316 6436 1324
rect 6492 1316 6500 1324
rect 4908 1296 4916 1304
rect 5948 1296 5956 1304
rect 6108 1296 6116 1304
rect 6172 1296 6180 1304
rect 6284 1296 6292 1304
rect 6572 1316 6580 1324
rect 6620 1316 6628 1324
rect 6668 1316 6676 1324
rect 6684 1316 6692 1324
rect 6716 1316 6724 1324
rect 6764 1316 6772 1324
rect 6780 1316 6788 1324
rect 6812 1316 6820 1324
rect 6892 1316 6900 1324
rect 7036 1316 7044 1324
rect 7228 1316 7236 1324
rect 6892 1296 6900 1304
rect 7308 1296 7316 1304
rect 588 1276 596 1284
rect 3564 1276 3572 1284
rect 3852 1276 3860 1284
rect 3964 1276 3972 1284
rect 4060 1276 4068 1284
rect 6076 1276 6084 1284
rect 6396 1276 6404 1284
rect 6524 1276 6532 1284
rect 6844 1276 6852 1284
rect 6924 1276 6932 1284
rect 604 1256 612 1264
rect 5116 1256 5124 1264
rect 188 1236 196 1244
rect 476 1236 484 1244
rect 1612 1236 1620 1244
rect 2828 1236 2836 1244
rect 3020 1236 3028 1244
rect 3276 1236 3284 1244
rect 3436 1236 3444 1244
rect 3484 1236 3492 1244
rect 3644 1236 3652 1244
rect 3692 1236 3700 1244
rect 3772 1236 3780 1244
rect 4204 1236 4212 1244
rect 5132 1236 5140 1244
rect 5180 1236 5188 1244
rect 5404 1236 5412 1244
rect 5468 1236 5476 1244
rect 5564 1236 5572 1244
rect 5644 1236 5652 1244
rect 5916 1236 5924 1244
rect 6572 1236 6580 1244
rect 7324 1236 7332 1244
rect 1411 1206 1419 1214
rect 1421 1206 1429 1214
rect 1431 1206 1439 1214
rect 1441 1206 1449 1214
rect 1451 1206 1459 1214
rect 1461 1206 1469 1214
rect 4419 1206 4427 1214
rect 4429 1206 4437 1214
rect 4439 1206 4447 1214
rect 4449 1206 4457 1214
rect 4459 1206 4467 1214
rect 4469 1206 4477 1214
rect 204 1176 212 1184
rect 268 1176 276 1184
rect 1020 1176 1028 1184
rect 1580 1176 1588 1184
rect 1756 1176 1764 1184
rect 1932 1176 1940 1184
rect 1948 1176 1956 1184
rect 2012 1176 2020 1184
rect 2076 1176 2084 1184
rect 2140 1176 2148 1184
rect 2204 1176 2212 1184
rect 2252 1176 2260 1184
rect 2300 1176 2308 1184
rect 2380 1176 2388 1184
rect 2396 1176 2404 1184
rect 2508 1176 2516 1184
rect 2524 1176 2532 1184
rect 2620 1176 2628 1184
rect 3564 1176 3572 1184
rect 3980 1176 3988 1184
rect 4012 1176 4020 1184
rect 4108 1176 4116 1184
rect 4220 1176 4228 1184
rect 4236 1176 4244 1184
rect 4300 1176 4308 1184
rect 4476 1176 4484 1184
rect 4540 1176 4548 1184
rect 4556 1176 4564 1184
rect 4620 1176 4628 1184
rect 4716 1176 4724 1184
rect 4796 1176 4804 1184
rect 4812 1176 4820 1184
rect 5084 1176 5092 1184
rect 5532 1176 5540 1184
rect 5628 1176 5636 1184
rect 5820 1176 5828 1184
rect 6012 1176 6020 1184
rect 6252 1176 6260 1184
rect 6268 1176 6276 1184
rect 6572 1176 6580 1184
rect 6764 1176 6772 1184
rect 4428 1156 4436 1164
rect 4684 1156 4692 1164
rect 6140 1156 6148 1164
rect 732 1136 740 1144
rect 1660 1136 1668 1144
rect 2572 1136 2580 1144
rect 4092 1136 4100 1144
rect 4252 1136 4260 1144
rect 4332 1136 4340 1144
rect 4588 1136 4596 1144
rect 4652 1136 4660 1144
rect 4732 1136 4740 1144
rect 4828 1136 4836 1144
rect 4860 1136 4868 1144
rect 5324 1136 5332 1144
rect 6972 1136 6980 1144
rect 7052 1136 7060 1144
rect 172 1116 180 1124
rect 668 1116 676 1124
rect 844 1116 852 1124
rect 940 1116 948 1124
rect 1148 1116 1156 1124
rect 1308 1116 1316 1124
rect 1740 1116 1748 1124
rect 1772 1116 1780 1124
rect 1852 1116 1860 1124
rect 2860 1116 2868 1124
rect 3436 1116 3444 1124
rect 3884 1116 3892 1124
rect 4028 1116 4036 1124
rect 4124 1116 4132 1124
rect 4172 1116 4180 1124
rect 4284 1116 4292 1124
rect 4348 1116 4356 1124
rect 4364 1116 4372 1124
rect 4604 1116 4612 1124
rect 4668 1116 4676 1124
rect 4764 1116 4772 1124
rect 4860 1116 4868 1124
rect 5500 1116 5508 1124
rect 220 1096 228 1104
rect 268 1096 276 1104
rect 316 1096 324 1104
rect 364 1096 372 1104
rect 476 1096 484 1104
rect 492 1096 500 1104
rect 556 1096 564 1104
rect 652 1096 660 1104
rect 684 1096 692 1104
rect 748 1096 756 1104
rect 828 1096 836 1104
rect 876 1096 884 1104
rect 956 1096 964 1104
rect 988 1096 996 1104
rect 1084 1096 1092 1104
rect 1164 1096 1172 1104
rect 1260 1096 1268 1104
rect 1340 1096 1348 1104
rect 1420 1096 1428 1104
rect 1436 1096 1444 1104
rect 1564 1096 1572 1104
rect 1580 1096 1588 1104
rect 1932 1096 1940 1104
rect 1980 1096 1988 1104
rect 2028 1096 2036 1104
rect 2044 1096 2052 1104
rect 2124 1096 2132 1104
rect 2236 1096 2244 1104
rect 2284 1096 2292 1104
rect 2332 1096 2340 1104
rect 2348 1096 2356 1104
rect 2460 1096 2468 1104
rect 2556 1096 2564 1104
rect 2604 1096 2612 1104
rect 2652 1096 2660 1104
rect 2796 1094 2804 1102
rect 2908 1096 2916 1104
rect 3116 1094 3124 1102
rect 3228 1096 3236 1104
rect 3340 1096 3348 1104
rect 3468 1096 3476 1104
rect 3548 1096 3556 1104
rect 3692 1094 3700 1102
rect 3788 1096 3796 1104
rect 3932 1096 3940 1104
rect 4108 1096 4116 1104
rect 4220 1096 4228 1104
rect 4268 1096 4276 1104
rect 4332 1096 4340 1104
rect 4380 1096 4388 1104
rect 4588 1096 4596 1104
rect 4652 1096 4660 1104
rect 4748 1096 4756 1104
rect 4844 1096 4852 1104
rect 4956 1094 4964 1102
rect 5132 1096 5140 1104
rect 5212 1096 5220 1104
rect 5260 1096 5268 1104
rect 5340 1096 5348 1104
rect 5404 1096 5412 1104
rect 5452 1096 5460 1104
rect 5532 1096 5540 1104
rect 5708 1116 5716 1124
rect 6092 1116 6100 1124
rect 5596 1096 5604 1104
rect 5628 1096 5636 1104
rect 5676 1096 5684 1104
rect 5708 1096 5716 1104
rect 5724 1096 5732 1104
rect 5788 1096 5796 1104
rect 5884 1096 5892 1104
rect 5980 1096 5988 1104
rect 6028 1096 6036 1104
rect 6044 1096 6052 1104
rect 6492 1116 6500 1124
rect 6140 1096 6148 1104
rect 6172 1096 6180 1104
rect 6220 1096 6228 1104
rect 6332 1096 6340 1104
rect 6364 1096 6372 1104
rect 7004 1116 7012 1124
rect 6524 1096 6532 1104
rect 6540 1096 6548 1104
rect 6636 1096 6644 1104
rect 6684 1096 6692 1104
rect 6828 1096 6836 1104
rect 6860 1096 6868 1104
rect 6972 1096 6980 1104
rect 7100 1096 7108 1104
rect 7116 1096 7124 1104
rect 7244 1096 7252 1104
rect 7308 1096 7316 1104
rect 7372 1096 7380 1104
rect 12 1076 20 1084
rect 60 1076 68 1084
rect 156 1076 164 1084
rect 220 1076 228 1084
rect 284 1076 292 1084
rect 428 1076 436 1084
rect 476 1076 484 1084
rect 508 1076 516 1084
rect 700 1076 708 1084
rect 860 1076 868 1084
rect 892 1076 900 1084
rect 908 1076 916 1084
rect 1020 1076 1028 1084
rect 1052 1076 1060 1084
rect 1116 1076 1124 1084
rect 236 1056 244 1064
rect 332 1056 340 1064
rect 380 1056 388 1064
rect 588 1056 596 1064
rect 636 1056 644 1064
rect 652 1056 660 1064
rect 732 1056 740 1064
rect 780 1056 788 1064
rect 988 1056 996 1064
rect 1084 1056 1092 1064
rect 1356 1076 1364 1084
rect 1372 1076 1380 1084
rect 1404 1076 1412 1084
rect 1516 1076 1524 1084
rect 1628 1076 1636 1084
rect 1724 1076 1732 1084
rect 1772 1076 1780 1084
rect 1820 1076 1828 1084
rect 1852 1076 1860 1084
rect 2172 1080 2180 1088
rect 2188 1076 2196 1084
rect 2428 1076 2436 1084
rect 2460 1076 2468 1084
rect 2876 1076 2884 1084
rect 2908 1076 2916 1084
rect 3212 1076 3220 1084
rect 3356 1076 3364 1084
rect 3452 1076 3460 1084
rect 3500 1076 3508 1084
rect 3532 1076 3540 1084
rect 3676 1076 3684 1084
rect 3916 1076 3924 1084
rect 3948 1076 3956 1084
rect 4060 1076 4068 1084
rect 4140 1076 4148 1084
rect 4924 1076 4932 1084
rect 5132 1076 5140 1084
rect 5356 1076 5364 1084
rect 5452 1076 5460 1084
rect 5516 1076 5524 1084
rect 5580 1076 5588 1084
rect 5644 1076 5652 1084
rect 5660 1076 5668 1084
rect 5724 1076 5732 1084
rect 5772 1076 5780 1084
rect 5836 1076 5844 1084
rect 6060 1076 6068 1084
rect 6156 1076 6164 1084
rect 6460 1076 6468 1084
rect 6556 1076 6564 1084
rect 6732 1076 6740 1084
rect 6956 1076 6964 1084
rect 7212 1076 7220 1084
rect 7260 1076 7268 1084
rect 7292 1076 7300 1084
rect 7356 1076 7364 1084
rect 1228 1056 1236 1064
rect 1276 1056 1284 1064
rect 1372 1056 1380 1064
rect 1516 1056 1524 1064
rect 1532 1056 1540 1064
rect 1612 1056 1620 1064
rect 1836 1056 1844 1064
rect 1852 1056 1860 1064
rect 1900 1056 1908 1064
rect 1996 1056 2004 1064
rect 2076 1056 2084 1064
rect 2444 1056 2452 1064
rect 2508 1056 2516 1064
rect 2524 1056 2532 1064
rect 2796 1056 2804 1064
rect 3116 1056 3124 1064
rect 3180 1056 3188 1064
rect 3500 1056 3508 1064
rect 3804 1056 3812 1064
rect 3868 1056 3876 1064
rect 3980 1056 3988 1064
rect 3996 1056 4004 1064
rect 4188 1056 4196 1064
rect 4508 1056 4516 1064
rect 4524 1056 4532 1064
rect 4700 1056 4708 1064
rect 4780 1056 4788 1064
rect 4892 1056 4900 1064
rect 5100 1056 5108 1064
rect 5132 1056 5140 1064
rect 5436 1056 5444 1064
rect 5756 1056 5764 1064
rect 5852 1056 5860 1064
rect 6204 1056 6212 1064
rect 7148 1056 7156 1064
rect 7212 1056 7220 1064
rect 7324 1056 7332 1064
rect 124 1036 132 1044
rect 460 1036 468 1044
rect 524 1036 532 1044
rect 796 1036 804 1044
rect 924 1036 932 1044
rect 972 1036 980 1044
rect 1100 1036 1108 1044
rect 1196 1036 1204 1044
rect 1292 1036 1300 1044
rect 1308 1036 1316 1044
rect 2092 1036 2100 1044
rect 2668 1036 2676 1044
rect 2924 1036 2932 1044
rect 3196 1036 3204 1044
rect 3244 1036 3252 1044
rect 3516 1036 3524 1044
rect 3564 1036 3572 1044
rect 3756 1036 3764 1044
rect 3852 1036 3860 1044
rect 3900 1036 3908 1044
rect 4044 1036 4052 1044
rect 5372 1036 5380 1044
rect 5500 1036 5508 1044
rect 6188 1036 6196 1044
rect 6252 1036 6260 1044
rect 6764 1036 6772 1044
rect 7020 1036 7028 1044
rect 7340 1036 7348 1044
rect 2915 1006 2923 1014
rect 2925 1006 2933 1014
rect 2935 1006 2943 1014
rect 2945 1006 2953 1014
rect 2955 1006 2963 1014
rect 2965 1006 2973 1014
rect 5923 1006 5931 1014
rect 5933 1006 5941 1014
rect 5943 1006 5951 1014
rect 5953 1006 5961 1014
rect 5963 1006 5971 1014
rect 5973 1006 5981 1014
rect 108 976 116 984
rect 236 976 244 984
rect 700 976 708 984
rect 796 976 804 984
rect 908 976 916 984
rect 1276 976 1284 984
rect 1388 976 1396 984
rect 1676 976 1684 984
rect 2012 976 2020 984
rect 2044 976 2052 984
rect 2188 976 2196 984
rect 2204 976 2212 984
rect 2284 976 2292 984
rect 2364 976 2372 984
rect 2460 976 2468 984
rect 2492 976 2500 984
rect 2620 976 2628 984
rect 2988 976 2996 984
rect 3228 976 3236 984
rect 3420 976 3428 984
rect 3500 976 3508 984
rect 3948 976 3956 984
rect 4236 976 4244 984
rect 4284 976 4292 984
rect 4620 976 4628 984
rect 4668 976 4676 984
rect 4940 976 4948 984
rect 5116 976 5124 984
rect 5676 976 5684 984
rect 5740 976 5748 984
rect 6236 976 6244 984
rect 6508 976 6516 984
rect 7004 976 7012 984
rect 7052 976 7060 984
rect 7324 976 7332 984
rect 396 956 404 964
rect 476 956 484 964
rect 524 956 532 964
rect 540 956 548 964
rect 572 956 580 964
rect 732 956 740 964
rect 764 956 772 964
rect 892 956 900 964
rect 956 956 964 964
rect 1116 956 1124 964
rect 1228 956 1236 964
rect 1740 956 1748 964
rect 1996 956 2004 964
rect 2108 956 2116 964
rect 2332 956 2340 964
rect 2428 956 2436 964
rect 2476 956 2484 964
rect 2636 956 2644 964
rect 3356 956 3364 964
rect 3484 956 3492 964
rect 3724 956 3732 964
rect 3932 956 3940 964
rect 3964 956 3972 964
rect 4044 956 4052 964
rect 4092 956 4100 964
rect 4124 956 4132 964
rect 4252 956 4260 964
rect 4652 956 4660 964
rect 4860 956 4868 964
rect 4924 956 4932 964
rect 5420 956 5428 964
rect 6140 956 6148 964
rect 6268 956 6276 964
rect 6604 956 6612 964
rect 6668 956 6676 964
rect 6764 956 6772 964
rect 7292 956 7300 964
rect 7340 956 7348 964
rect 60 936 68 944
rect 156 936 164 944
rect 172 936 180 944
rect 268 936 276 944
rect 284 936 292 944
rect 364 936 372 944
rect 620 936 628 944
rect 652 936 660 944
rect 716 936 724 944
rect 812 936 820 944
rect 924 936 932 944
rect 940 936 948 944
rect 1036 936 1044 944
rect 1052 936 1060 944
rect 1068 936 1076 944
rect 1324 936 1332 944
rect 1340 936 1348 944
rect 1436 936 1444 944
rect 1516 936 1524 944
rect 1628 936 1636 944
rect 1724 936 1732 944
rect 1820 936 1828 944
rect 1932 936 1940 944
rect 2076 932 2084 940
rect 2092 936 2100 944
rect 2140 936 2148 944
rect 2268 936 2276 944
rect 2796 936 2804 944
rect 2844 936 2852 944
rect 3116 936 3124 944
rect 3196 936 3204 944
rect 3388 936 3396 944
rect 3468 936 3476 944
rect 3516 936 3524 944
rect 3596 936 3604 944
rect 3692 936 3700 944
rect 3836 936 3844 944
rect 3900 936 3908 944
rect 3932 936 3940 944
rect 3996 936 4004 944
rect 4172 936 4180 944
rect 4188 936 4196 944
rect 4444 936 4452 944
rect 4540 936 4548 944
rect 4604 936 4612 944
rect 4684 936 4692 944
rect 4748 936 4756 944
rect 4796 936 4804 944
rect 4860 936 4868 944
rect 4892 936 4900 944
rect 4956 936 4964 944
rect 5020 936 5028 944
rect 5068 936 5076 944
rect 5180 936 5188 944
rect 5212 936 5220 944
rect 5244 936 5252 944
rect 5276 936 5284 944
rect 5308 936 5316 944
rect 5468 936 5476 944
rect 5532 936 5540 944
rect 5548 936 5556 944
rect 5868 936 5876 944
rect 5980 936 5988 944
rect 6124 936 6132 944
rect 6188 936 6196 944
rect 6252 936 6260 944
rect 6332 936 6340 944
rect 6428 936 6436 944
rect 6476 936 6484 944
rect 6492 936 6500 944
rect 6556 936 6564 944
rect 6620 936 6628 944
rect 6684 936 6692 944
rect 6748 936 6756 944
rect 7036 936 7044 944
rect 7148 936 7156 944
rect 7244 936 7252 944
rect 7308 936 7316 944
rect 44 916 52 924
rect 316 916 324 924
rect 444 916 452 924
rect 492 916 500 924
rect 572 916 580 924
rect 636 916 644 924
rect 668 916 676 924
rect 332 896 340 904
rect 732 916 740 924
rect 860 916 868 924
rect 956 916 964 924
rect 1020 916 1028 924
rect 1164 916 1172 924
rect 1212 916 1220 924
rect 1260 916 1268 924
rect 1308 916 1316 924
rect 1756 916 1764 924
rect 1980 916 1988 924
rect 2028 916 2036 924
rect 2156 916 2164 924
rect 2236 916 2244 924
rect 2252 916 2260 924
rect 2380 916 2388 924
rect 2444 916 2452 924
rect 2524 916 2532 924
rect 2540 916 2548 924
rect 2588 916 2596 924
rect 2668 916 2676 924
rect 2812 918 2820 926
rect 2876 916 2884 924
rect 3020 916 3028 924
rect 3164 918 3172 926
rect 3356 918 3364 926
rect 3452 916 3460 924
rect 3532 916 3540 924
rect 3548 916 3556 924
rect 3612 916 3620 924
rect 3724 916 3732 924
rect 3772 916 3780 924
rect 3820 916 3828 924
rect 3884 916 3892 924
rect 3900 916 3908 924
rect 4012 916 4020 924
rect 4092 916 4100 924
rect 4124 916 4132 924
rect 4204 916 4212 924
rect 4348 916 4356 924
rect 4412 918 4420 926
rect 4844 916 4852 924
rect 4908 916 4916 924
rect 5020 916 5028 924
rect 5100 916 5108 924
rect 5148 916 5156 924
rect 5164 916 5172 924
rect 5180 916 5188 924
rect 5228 916 5236 924
rect 780 896 788 904
rect 876 896 884 904
rect 1004 896 1012 904
rect 1276 896 1284 904
rect 1788 896 1796 904
rect 3420 896 3428 904
rect 3644 896 3652 904
rect 3756 896 3764 904
rect 3868 896 3876 904
rect 3964 896 3972 904
rect 4140 896 4148 904
rect 4236 896 4244 904
rect 4572 896 4580 904
rect 4716 896 4724 904
rect 4748 896 4756 904
rect 4844 896 4852 904
rect 4988 896 4996 904
rect 5036 896 5044 904
rect 5308 916 5316 924
rect 5340 916 5348 924
rect 5388 916 5396 924
rect 5404 916 5412 924
rect 5452 916 5460 924
rect 5468 916 5476 924
rect 5516 916 5524 924
rect 5564 916 5572 924
rect 5612 916 5620 924
rect 5628 916 5636 924
rect 5660 916 5668 924
rect 5708 916 5716 924
rect 5724 916 5732 924
rect 5852 916 5860 924
rect 5996 916 6004 924
rect 6076 916 6084 924
rect 6108 916 6116 924
rect 6172 916 6180 924
rect 6188 916 6196 924
rect 6236 916 6244 924
rect 6300 916 6308 924
rect 6316 916 6324 924
rect 6396 916 6404 924
rect 6412 916 6420 924
rect 6444 916 6452 924
rect 6508 916 6516 924
rect 6556 916 6564 924
rect 6572 916 6580 924
rect 6620 916 6628 924
rect 5484 896 5492 904
rect 6044 896 6052 904
rect 6268 896 6276 904
rect 6476 896 6484 904
rect 6700 916 6708 924
rect 6796 916 6804 924
rect 6812 916 6820 924
rect 6828 916 6836 924
rect 6892 916 6900 924
rect 6908 916 6916 924
rect 6924 916 6932 924
rect 6988 916 6996 924
rect 7164 916 7172 924
rect 7244 916 7252 924
rect 7308 916 7316 924
rect 7004 896 7012 904
rect 12 876 20 884
rect 364 876 372 884
rect 396 876 404 884
rect 844 876 852 884
rect 1548 876 1556 884
rect 1868 876 1876 884
rect 2684 876 2692 884
rect 3036 876 3044 884
rect 3260 876 3268 884
rect 3788 876 3796 884
rect 4124 876 4132 884
rect 4764 876 4772 884
rect 4796 876 4804 884
rect 5452 876 5460 884
rect 6076 876 6084 884
rect 6172 876 6180 884
rect 6572 876 6580 884
rect 6668 876 6676 884
rect 860 856 868 864
rect 348 836 356 844
rect 460 836 468 844
rect 1132 836 1140 844
rect 1180 836 1188 844
rect 1228 836 1236 844
rect 1948 836 1956 844
rect 2124 836 2132 844
rect 2492 836 2500 844
rect 2572 836 2580 844
rect 2620 836 2628 844
rect 2908 836 2916 844
rect 3580 836 3588 844
rect 3660 836 3668 844
rect 3804 836 3812 844
rect 3948 836 3956 844
rect 4268 836 4276 844
rect 5356 836 5364 844
rect 6364 836 6372 844
rect 6700 836 6708 844
rect 6844 836 6852 844
rect 6940 836 6948 844
rect 1411 806 1419 814
rect 1421 806 1429 814
rect 1431 806 1439 814
rect 1441 806 1449 814
rect 1451 806 1459 814
rect 1461 806 1469 814
rect 4419 806 4427 814
rect 4429 806 4437 814
rect 4439 806 4447 814
rect 4449 806 4457 814
rect 4459 806 4467 814
rect 4469 806 4477 814
rect 12 776 20 784
rect 236 776 244 784
rect 940 776 948 784
rect 1020 776 1028 784
rect 1164 776 1172 784
rect 1276 776 1284 784
rect 1388 776 1396 784
rect 1900 776 1908 784
rect 2316 776 2324 784
rect 2412 776 2420 784
rect 2748 776 2756 784
rect 3196 776 3204 784
rect 3516 776 3524 784
rect 3852 776 3860 784
rect 4012 776 4020 784
rect 4060 776 4068 784
rect 4252 776 4260 784
rect 4316 776 4324 784
rect 4348 776 4356 784
rect 4508 776 4516 784
rect 4860 776 4868 784
rect 4892 776 4900 784
rect 5196 776 5204 784
rect 5516 776 5524 784
rect 5532 776 5540 784
rect 6220 776 6228 784
rect 6316 776 6324 784
rect 6604 776 6612 784
rect 6796 776 6804 784
rect 6988 776 6996 784
rect 7228 776 7236 784
rect 7356 776 7364 784
rect 2396 756 2404 764
rect 2476 756 2484 764
rect 2924 756 2932 764
rect 5820 756 5828 764
rect 6700 756 6708 764
rect 140 736 148 744
rect 284 736 292 744
rect 316 736 324 744
rect 572 736 580 744
rect 2492 736 2500 744
rect 2828 736 2836 744
rect 3020 736 3028 744
rect 3980 736 3988 744
rect 4156 736 4164 744
rect 4220 736 4228 744
rect 4716 736 4724 744
rect 4812 736 4820 744
rect 6124 736 6132 744
rect 6172 736 6180 744
rect 108 716 116 724
rect 172 716 180 724
rect 348 716 356 724
rect 460 716 468 724
rect 524 716 532 724
rect 540 716 548 724
rect 876 716 884 724
rect 1036 716 1044 724
rect 1292 716 1300 724
rect 1500 716 1508 724
rect 1532 716 1540 724
rect 1772 716 1780 724
rect 2188 716 2196 724
rect 2460 716 2468 724
rect 2572 716 2580 724
rect 2716 716 2724 724
rect 2780 716 2788 724
rect 3004 716 3012 724
rect 3068 716 3076 724
rect 3436 716 3444 724
rect 3756 716 3764 724
rect 3868 716 3876 724
rect 4044 716 4052 724
rect 4076 716 4084 724
rect 4124 716 4132 724
rect 4284 716 4292 724
rect 4732 716 4740 724
rect 4748 716 4756 724
rect 4844 716 4852 724
rect 5116 716 5124 724
rect 5292 716 5300 724
rect 5612 716 5620 724
rect 6412 716 6420 724
rect 6524 716 6532 724
rect 6908 716 6916 724
rect 7260 716 7268 724
rect 60 696 68 704
rect 156 696 164 704
rect 188 696 196 704
rect 284 696 292 704
rect 300 696 308 704
rect 364 696 372 704
rect 412 696 420 704
rect 476 696 484 704
rect 540 696 548 704
rect 572 696 580 704
rect 668 696 676 704
rect 764 696 772 704
rect 844 696 852 704
rect 876 696 884 704
rect 956 696 964 704
rect 1004 696 1012 704
rect 1244 696 1252 704
rect 1340 696 1348 704
rect 1516 696 1524 704
rect 1596 696 1604 704
rect 1612 696 1620 704
rect 1996 696 2004 704
rect 2140 696 2148 704
rect 2188 696 2196 704
rect 2236 696 2244 704
rect 2268 696 2276 704
rect 2284 696 2292 704
rect 2364 696 2372 704
rect 2412 696 2420 704
rect 2476 696 2484 704
rect 2556 696 2564 704
rect 2668 696 2676 704
rect 2748 696 2756 704
rect 2876 696 2884 704
rect 3052 696 3060 704
rect 3100 696 3108 704
rect 3180 696 3188 704
rect 3260 696 3268 704
rect 3324 694 3332 702
rect 3404 696 3412 704
rect 3500 696 3508 704
rect 3644 694 3652 702
rect 3724 696 3732 704
rect 3820 696 3828 704
rect 3900 696 3908 704
rect 3932 696 3940 704
rect 3996 696 4004 704
rect 4156 696 4164 704
rect 4236 696 4244 704
rect 4252 696 4260 704
rect 4636 694 4644 702
rect 4796 696 4804 704
rect 5020 694 5028 702
rect 5164 696 5172 704
rect 5244 696 5252 704
rect 5388 694 5396 702
rect 5452 696 5460 704
rect 5564 696 5572 704
rect 5708 694 5716 702
rect 5772 696 5780 704
rect 5836 696 5844 704
rect 6012 696 6020 704
rect 6140 696 6148 704
rect 6188 696 6196 704
rect 6204 696 6212 704
rect 6252 696 6260 704
rect 6300 696 6308 704
rect 6396 696 6404 704
rect 6444 696 6452 704
rect 6492 696 6500 704
rect 6556 696 6564 704
rect 6572 696 6580 704
rect 6604 696 6612 704
rect 6636 696 6644 704
rect 6684 696 6692 704
rect 6732 696 6740 704
rect 6748 696 6756 704
rect 6780 696 6788 704
rect 6828 696 6836 704
rect 6844 696 6852 704
rect 6860 696 6868 704
rect 6876 696 6884 704
rect 6924 696 6932 704
rect 6956 696 6964 704
rect 6972 696 6980 704
rect 7020 696 7028 704
rect 7052 696 7060 704
rect 7100 696 7108 704
rect 7148 696 7156 704
rect 7212 696 7220 704
rect 7228 696 7236 704
rect 7260 696 7268 704
rect 7324 696 7332 704
rect 7372 696 7380 704
rect 76 676 84 684
rect 156 676 164 684
rect 204 676 212 684
rect 300 676 308 684
rect 12 656 20 664
rect 236 656 244 664
rect 252 656 260 664
rect 364 656 372 664
rect 428 676 436 684
rect 460 676 468 684
rect 492 676 500 684
rect 588 676 596 684
rect 700 676 708 684
rect 716 676 724 684
rect 796 676 804 684
rect 844 676 852 684
rect 940 676 948 684
rect 1084 676 1092 684
rect 668 656 676 664
rect 780 656 788 664
rect 972 656 980 664
rect 1036 656 1044 664
rect 1116 676 1124 684
rect 1212 676 1220 684
rect 1228 676 1236 684
rect 1340 676 1348 684
rect 1356 676 1364 684
rect 1468 676 1476 684
rect 1388 656 1396 664
rect 1564 656 1572 664
rect 1580 656 1588 664
rect 1628 656 1636 664
rect 1740 676 1748 684
rect 1836 676 1844 684
rect 1852 676 1860 684
rect 1948 676 1956 684
rect 1996 676 2004 684
rect 2092 676 2100 684
rect 2156 676 2164 684
rect 2220 676 2228 684
rect 2252 676 2260 684
rect 2332 676 2340 684
rect 2620 676 2628 684
rect 2892 676 2900 684
rect 3036 676 3044 684
rect 3148 676 3156 684
rect 3388 676 3396 684
rect 3484 676 3492 684
rect 3676 676 3684 684
rect 3708 676 3716 684
rect 3804 676 3812 684
rect 3916 676 3924 684
rect 3948 676 3956 684
rect 4172 676 4180 684
rect 4220 676 4228 684
rect 4364 676 4372 684
rect 4540 676 4548 684
rect 4700 676 4708 684
rect 4780 676 4788 684
rect 4812 676 4820 684
rect 4924 676 4932 684
rect 5084 676 5092 684
rect 5148 676 5156 684
rect 5260 676 5268 684
rect 5324 676 5332 684
rect 5644 676 5652 684
rect 5740 676 5748 684
rect 5788 676 5796 684
rect 5868 676 5876 684
rect 6012 676 6020 684
rect 6268 676 6276 684
rect 6364 676 6372 684
rect 6396 676 6404 684
rect 6476 676 6484 684
rect 6540 676 6548 684
rect 6588 676 6596 684
rect 6668 676 6676 684
rect 7068 676 7076 684
rect 1660 656 1668 664
rect 1724 656 1732 664
rect 1980 656 1988 664
rect 2380 656 2388 664
rect 2444 656 2452 664
rect 2524 656 2532 664
rect 2636 656 2644 664
rect 2796 656 2804 664
rect 2828 656 2836 664
rect 2860 656 2868 664
rect 2940 656 2948 664
rect 3084 656 3092 664
rect 3228 656 3236 664
rect 3836 656 3844 664
rect 3980 656 3988 664
rect 4076 656 4084 664
rect 4108 656 4116 664
rect 4188 656 4196 664
rect 4300 656 4308 664
rect 4332 656 4340 664
rect 4636 656 4644 664
rect 4748 656 4756 664
rect 4844 656 4852 664
rect 4876 656 4884 664
rect 5020 656 5028 664
rect 5180 656 5188 664
rect 5212 656 5220 664
rect 5228 656 5236 664
rect 5932 656 5940 664
rect 6364 656 6372 664
rect 6540 656 6548 664
rect 7212 676 7220 684
rect 7308 676 7316 684
rect 7116 656 7124 664
rect 7148 656 7156 664
rect 7196 656 7204 664
rect 7276 656 7284 664
rect 7340 656 7348 664
rect 108 636 116 644
rect 684 636 692 644
rect 1292 636 1300 644
rect 1484 636 1492 644
rect 1676 636 1684 644
rect 1964 636 1972 644
rect 2108 636 2116 644
rect 2188 636 2196 644
rect 3132 636 3140 644
rect 3468 636 3476 644
rect 3788 636 3796 644
rect 3868 636 3876 644
rect 4380 636 4388 644
rect 5580 636 5588 644
rect 2915 606 2923 614
rect 2925 606 2933 614
rect 2935 606 2943 614
rect 2945 606 2953 614
rect 2955 606 2963 614
rect 2965 606 2973 614
rect 5923 606 5931 614
rect 5933 606 5941 614
rect 5943 606 5951 614
rect 5953 606 5961 614
rect 5963 606 5971 614
rect 5973 606 5981 614
rect 156 576 164 584
rect 572 576 580 584
rect 844 576 852 584
rect 1020 576 1028 584
rect 1100 576 1108 584
rect 1356 576 1364 584
rect 1564 576 1572 584
rect 1788 576 1796 584
rect 2204 576 2212 584
rect 2460 576 2468 584
rect 2748 576 2756 584
rect 2892 576 2900 584
rect 3164 576 3172 584
rect 3612 576 3620 584
rect 4204 576 4212 584
rect 4220 576 4228 584
rect 4524 576 4532 584
rect 4796 576 4804 584
rect 4924 576 4932 584
rect 5484 576 5492 584
rect 5740 576 5748 584
rect 6140 576 6148 584
rect 6156 576 6164 584
rect 6748 576 6756 584
rect 6924 576 6932 584
rect 7180 576 7188 584
rect 12 556 20 564
rect 44 556 52 564
rect 60 556 68 564
rect 76 556 84 564
rect 364 556 372 564
rect 380 556 388 564
rect 444 556 452 564
rect 556 556 564 564
rect 668 556 676 564
rect 684 556 692 564
rect 700 556 708 564
rect 780 556 788 564
rect 988 556 996 564
rect 1004 556 1012 564
rect 1180 556 1188 564
rect 1212 556 1220 564
rect 1644 556 1652 564
rect 1708 556 1716 564
rect 1772 556 1780 564
rect 1836 556 1844 564
rect 1948 556 1956 564
rect 2092 556 2100 564
rect 2188 556 2196 564
rect 2252 556 2260 564
rect 2364 556 2372 564
rect 2428 556 2436 564
rect 2588 556 2596 564
rect 2876 556 2884 564
rect 2908 556 2916 564
rect 3036 556 3044 564
rect 3820 556 3828 564
rect 3836 556 3844 564
rect 3900 556 3908 564
rect 3980 556 3988 564
rect 4812 556 4820 564
rect 4876 556 4884 564
rect 5212 556 5220 564
rect 5308 556 5316 564
rect 5468 556 5476 564
rect 5676 556 5684 564
rect 5788 556 5796 564
rect 6012 556 6020 564
rect 6620 556 6628 564
rect 188 536 196 544
rect 252 536 260 544
rect 284 536 292 544
rect 412 536 420 544
rect 588 536 596 544
rect 620 536 628 544
rect 700 536 708 544
rect 748 536 756 544
rect 796 536 804 544
rect 860 536 868 544
rect 908 536 916 544
rect 1036 536 1044 544
rect 12 516 20 524
rect 44 516 52 524
rect 236 516 244 524
rect 268 516 276 524
rect 300 516 308 524
rect 332 516 340 524
rect 492 516 500 524
rect 540 516 548 524
rect 1164 536 1172 544
rect 1260 536 1268 544
rect 1292 536 1300 544
rect 1340 536 1348 544
rect 1420 536 1428 544
rect 1516 536 1524 544
rect 1532 536 1540 544
rect 1628 536 1636 544
rect 1676 536 1684 544
rect 1708 536 1716 544
rect 1868 536 1876 544
rect 1980 536 1988 544
rect 2012 536 2020 544
rect 2028 536 2036 544
rect 2108 536 2116 544
rect 2140 536 2148 544
rect 2188 536 2196 544
rect 2364 536 2372 544
rect 2396 536 2404 544
rect 2444 536 2452 544
rect 2492 536 2500 544
rect 2556 536 2564 544
rect 2652 536 2660 544
rect 2780 536 2788 544
rect 2812 536 2820 544
rect 2844 536 2852 544
rect 3020 536 3028 544
rect 3052 536 3060 544
rect 3260 536 3268 544
rect 3708 536 3716 544
rect 3964 536 3972 544
rect 4636 536 4644 544
rect 4684 536 4692 544
rect 4716 536 4724 544
rect 4780 536 4788 544
rect 4860 536 4868 544
rect 5020 536 5028 544
rect 5116 536 5124 544
rect 5180 536 5188 544
rect 5212 536 5220 544
rect 5372 536 5380 544
rect 5404 536 5412 544
rect 5436 536 5444 544
rect 5580 536 5588 544
rect 5644 536 5652 544
rect 5788 536 5796 544
rect 5820 536 5828 544
rect 5948 536 5956 544
rect 6348 536 6356 544
rect 6380 536 6388 544
rect 6444 536 6452 544
rect 6460 536 6468 544
rect 6556 536 6564 544
rect 6796 536 6804 544
rect 6812 536 6820 544
rect 6908 536 6916 544
rect 7052 536 7060 544
rect 7116 536 7124 544
rect 7148 536 7156 544
rect 668 516 676 524
rect 844 516 852 524
rect 876 516 884 524
rect 956 516 964 524
rect 1052 516 1060 524
rect 1228 516 1236 524
rect 1276 516 1284 524
rect 1324 516 1332 524
rect 1388 516 1396 524
rect 1404 516 1412 524
rect 1500 516 1508 524
rect 1596 516 1604 524
rect 1692 516 1700 524
rect 1820 516 1828 524
rect 1916 516 1924 524
rect 2060 516 2068 524
rect 2156 516 2164 524
rect 2220 516 2228 524
rect 2236 516 2244 524
rect 2300 516 2308 524
rect 2316 516 2324 524
rect 2508 516 2516 524
rect 2524 516 2532 524
rect 2540 516 2548 524
rect 2636 516 2644 524
rect 2684 516 2692 524
rect 2732 516 2740 524
rect 2796 516 2804 524
rect 3148 516 3156 524
rect 3292 518 3300 526
rect 3420 516 3428 524
rect 3484 518 3492 526
rect 3580 516 3588 524
rect 3740 518 3748 526
rect 3804 516 3812 524
rect 3868 516 3876 524
rect 3932 516 3940 524
rect 3948 516 3956 524
rect 4012 516 4020 524
rect 4076 518 4084 526
rect 4140 516 4148 524
rect 4284 516 4292 524
rect 4316 516 4324 524
rect 4412 516 4420 524
rect 4652 518 4660 526
rect 4908 516 4916 524
rect 5052 518 5060 526
rect 5196 516 5204 524
rect 5260 516 5268 524
rect 5276 516 5284 524
rect 5324 516 5332 524
rect 5468 516 5476 524
rect 5596 516 5604 524
rect 5708 516 5716 524
rect 5772 516 5780 524
rect 5804 516 5812 524
rect 6012 518 6020 526
rect 6076 516 6084 524
rect 6220 516 6228 524
rect 6284 518 6292 526
rect 204 496 212 504
rect 380 496 388 504
rect 412 496 420 504
rect 652 496 660 504
rect 716 496 724 504
rect 748 496 756 504
rect 876 496 884 504
rect 972 496 980 504
rect 1308 496 1316 504
rect 1420 496 1428 504
rect 1468 496 1476 504
rect 2396 496 2404 504
rect 2428 496 2436 504
rect 2476 496 2484 504
rect 2748 496 2756 504
rect 2812 496 2820 504
rect 3916 496 3924 504
rect 4748 496 4756 504
rect 4828 496 4836 504
rect 4844 496 4852 504
rect 5148 496 5156 504
rect 5372 496 5380 504
rect 5852 496 5860 504
rect 6380 496 6388 504
rect 6428 516 6436 524
rect 6492 496 6500 504
rect 6524 516 6532 524
rect 6556 516 6564 524
rect 6620 518 6628 526
rect 6684 516 6692 524
rect 6764 496 6772 504
rect 6844 496 6852 504
rect 6892 516 6900 524
rect 7036 516 7044 524
rect 7132 516 7140 524
rect 7244 516 7252 524
rect 7292 516 7300 524
rect 6892 496 6900 504
rect 7164 496 7172 504
rect 236 476 244 484
rect 2252 476 2260 484
rect 4012 476 4020 484
rect 460 436 468 444
rect 508 436 516 444
rect 924 436 932 444
rect 1196 436 1204 444
rect 1852 436 1860 444
rect 1916 436 1924 444
rect 2604 436 2612 444
rect 2700 436 2708 444
rect 3116 436 3124 444
rect 3356 436 3364 444
rect 3548 436 3556 444
rect 3868 436 3876 444
rect 4508 436 4516 444
rect 6780 436 6788 444
rect 1411 406 1419 414
rect 1421 406 1429 414
rect 1431 406 1439 414
rect 1441 406 1449 414
rect 1451 406 1459 414
rect 1461 406 1469 414
rect 4419 406 4427 414
rect 4429 406 4437 414
rect 4439 406 4447 414
rect 4449 406 4457 414
rect 4459 406 4467 414
rect 4469 406 4477 414
rect 44 376 52 384
rect 140 376 148 384
rect 1068 376 1076 384
rect 1084 376 1092 384
rect 1324 376 1332 384
rect 1356 376 1364 384
rect 1644 376 1652 384
rect 1756 376 1764 384
rect 2156 376 2164 384
rect 2236 376 2244 384
rect 2268 376 2276 384
rect 2492 376 2500 384
rect 3772 376 3780 384
rect 3916 376 3924 384
rect 4108 376 4116 384
rect 4220 376 4228 384
rect 4716 376 4724 384
rect 4812 376 4820 384
rect 4860 376 4868 384
rect 4972 376 4980 384
rect 5020 376 5028 384
rect 5244 376 5252 384
rect 5500 376 5508 384
rect 5900 376 5908 384
rect 6204 376 6212 384
rect 6252 376 6260 384
rect 6956 376 6964 384
rect 7004 376 7012 384
rect 7356 376 7364 384
rect 1612 356 1620 364
rect 2620 356 2628 364
rect 4476 356 4484 364
rect 844 336 852 344
rect 956 336 964 344
rect 1260 336 1268 344
rect 1868 336 1876 344
rect 2508 336 2516 344
rect 3340 336 3348 344
rect 3404 336 3412 344
rect 4796 336 4804 344
rect 5148 336 5156 344
rect 5420 336 5428 344
rect 6556 336 6564 344
rect 6732 336 6740 344
rect 188 316 196 324
rect 220 316 228 324
rect 364 316 372 324
rect 572 316 580 324
rect 796 316 804 324
rect 812 316 820 324
rect 892 316 900 324
rect 924 316 932 324
rect 1004 316 1012 324
rect 1148 316 1156 324
rect 1180 316 1188 324
rect 1276 316 1284 324
rect 1596 316 1604 324
rect 1628 316 1636 324
rect 1692 316 1700 324
rect 1836 316 1844 324
rect 1932 316 1940 324
rect 2220 316 2228 324
rect 2364 316 2372 324
rect 2476 316 2484 324
rect 2732 316 2740 324
rect 2876 316 2884 324
rect 3004 316 3012 324
rect 3068 316 3076 324
rect 3100 316 3108 324
rect 3884 316 3892 324
rect 3996 316 4004 324
rect 4044 316 4052 324
rect 4124 316 4132 324
rect 4172 316 4180 324
rect 4700 316 4708 324
rect 4908 316 4916 324
rect 5436 316 5444 324
rect 5596 316 5604 324
rect 5740 316 5748 324
rect 5788 316 5796 324
rect 5836 316 5844 324
rect 140 296 148 304
rect 236 296 244 304
rect 268 296 276 304
rect 300 296 308 304
rect 396 296 404 304
rect 428 296 436 304
rect 540 296 548 304
rect 572 296 580 304
rect 684 296 692 304
rect 764 296 772 304
rect 844 296 852 304
rect 956 296 964 304
rect 988 296 996 304
rect 1020 296 1028 304
rect 1132 296 1140 304
rect 1180 296 1188 304
rect 1324 296 1332 304
rect 1404 296 1412 304
rect 1548 296 1556 304
rect 1580 296 1588 304
rect 1788 296 1796 304
rect 1836 296 1844 304
rect 1916 296 1924 304
rect 2012 296 2020 304
rect 2204 296 2212 304
rect 2300 296 2308 304
rect 2348 296 2356 304
rect 2364 296 2372 304
rect 2412 296 2420 304
rect 2460 296 2468 304
rect 2492 296 2500 304
rect 2636 296 2644 304
rect 2716 296 2724 304
rect 2844 296 2852 304
rect 2908 296 2916 304
rect 2924 296 2932 304
rect 3052 296 3060 304
rect 3116 296 3124 304
rect 3148 296 3156 304
rect 3228 296 3236 304
rect 3292 296 3300 304
rect 12 276 20 284
rect 108 276 116 284
rect 124 276 132 284
rect 188 276 196 284
rect 204 276 212 284
rect 220 276 228 284
rect 3532 294 3540 302
rect 3660 296 3668 304
rect 3708 296 3716 304
rect 3788 296 3796 304
rect 3932 296 3940 304
rect 4284 296 4292 304
rect 4332 296 4340 304
rect 4588 296 4596 304
rect 4700 296 4708 304
rect 4748 296 4756 304
rect 4956 296 4964 304
rect 5276 296 5284 304
rect 5372 296 5380 304
rect 5388 296 5396 304
rect 5660 296 5668 304
rect 5740 296 5748 304
rect 5772 296 5780 304
rect 6092 296 6100 304
rect 6140 296 6148 304
rect 6284 296 6292 304
rect 6332 316 6340 324
rect 6764 316 6772 324
rect 6972 316 6980 324
rect 6428 294 6436 302
rect 6476 296 6484 304
rect 6572 296 6580 304
rect 6732 296 6740 304
rect 6828 294 6836 302
rect 7004 296 7012 304
rect 7260 296 7268 304
rect 476 276 484 284
rect 508 276 516 284
rect 588 276 596 284
rect 604 276 612 284
rect 636 276 644 284
rect 716 276 724 284
rect 860 276 868 284
rect 972 276 980 284
rect 1116 276 1124 284
rect 1196 276 1204 284
rect 1228 276 1236 284
rect 1244 276 1252 284
rect 1532 276 1540 284
rect 1596 276 1604 284
rect 1708 276 1716 284
rect 1772 276 1780 284
rect 1852 276 1860 284
rect 1868 276 1876 284
rect 1964 276 1972 284
rect 2028 276 2036 284
rect 2124 276 2132 284
rect 2172 276 2180 284
rect 2252 276 2260 284
rect 2412 276 2420 284
rect 2428 276 2436 284
rect 2540 276 2548 284
rect 2588 276 2596 284
rect 2764 276 2772 284
rect 2956 276 2964 284
rect 3068 276 3076 284
rect 3228 276 3236 284
rect 3276 276 3284 284
rect 3340 276 3348 284
rect 3484 276 3492 284
rect 3788 276 3796 284
rect 3852 276 3860 284
rect 3964 276 3972 284
rect 4028 276 4036 284
rect 4076 276 4084 284
rect 4156 276 4164 284
rect 4204 276 4212 284
rect 4380 276 4388 284
rect 4540 276 4548 284
rect 4636 276 4644 284
rect 4668 276 4676 284
rect 4732 276 4740 284
rect 4876 276 4884 284
rect 5132 276 5140 284
rect 5196 276 5204 284
rect 5356 276 5364 284
rect 5468 276 5476 284
rect 5548 276 5556 284
rect 5612 276 5620 284
rect 5708 276 5716 284
rect 5788 276 5796 284
rect 5820 276 5828 284
rect 5868 276 5876 284
rect 5884 276 5892 284
rect 6076 276 6084 284
rect 6268 276 6276 284
rect 6332 276 6340 284
rect 6364 276 6372 284
rect 6700 276 6708 284
rect 6716 276 6724 284
rect 6860 276 6868 284
rect 7020 276 7028 284
rect 7036 276 7044 284
rect 7164 276 7172 284
rect 7196 276 7204 284
rect 7244 276 7252 284
rect 332 256 340 264
rect 348 256 356 264
rect 396 256 404 264
rect 668 256 676 264
rect 716 256 724 264
rect 780 256 788 264
rect 908 256 916 264
rect 1020 256 1028 264
rect 1084 256 1092 264
rect 1212 256 1220 264
rect 1292 256 1300 264
rect 1420 256 1428 264
rect 1660 256 1668 264
rect 1980 256 1988 264
rect 2140 256 2148 264
rect 2540 256 2548 264
rect 2668 256 2676 264
rect 2796 256 2804 264
rect 3116 256 3124 264
rect 3148 256 3156 264
rect 3164 256 3172 264
rect 3372 256 3380 264
rect 3836 256 3844 264
rect 3868 256 3876 264
rect 3900 256 3908 264
rect 3932 256 3940 264
rect 4044 256 4052 264
rect 4092 256 4100 264
rect 4732 256 4740 264
rect 4796 256 4804 264
rect 4828 256 4836 264
rect 4844 256 4852 264
rect 4924 256 4932 264
rect 4988 256 4996 264
rect 5340 256 5348 264
rect 5436 256 5444 264
rect 5660 256 5668 264
rect 380 236 388 244
rect 428 236 436 244
rect 620 236 628 244
rect 732 236 740 244
rect 1612 236 1620 244
rect 1996 236 2004 244
rect 2092 236 2100 244
rect 2316 236 2324 244
rect 3196 236 3204 244
rect 3820 236 3828 244
rect 4124 236 4132 244
rect 4172 236 4180 244
rect 4908 236 4916 244
rect 5308 236 5316 244
rect 5692 236 5700 244
rect 5740 236 5748 244
rect 5836 236 5844 244
rect 2915 206 2923 214
rect 2925 206 2933 214
rect 2935 206 2943 214
rect 2945 206 2953 214
rect 2955 206 2963 214
rect 2965 206 2973 214
rect 5923 206 5931 214
rect 5933 206 5941 214
rect 5943 206 5951 214
rect 5953 206 5961 214
rect 5963 206 5971 214
rect 5973 206 5981 214
rect 60 176 68 184
rect 124 176 132 184
rect 188 176 196 184
rect 220 176 228 184
rect 284 176 292 184
rect 460 176 468 184
rect 636 176 644 184
rect 668 176 676 184
rect 764 176 772 184
rect 892 176 900 184
rect 1164 176 1172 184
rect 1260 176 1268 184
rect 1340 176 1348 184
rect 1644 176 1652 184
rect 1772 176 1780 184
rect 1836 176 1844 184
rect 2028 176 2036 184
rect 2108 176 2116 184
rect 2316 176 2324 184
rect 2348 176 2356 184
rect 2460 176 2468 184
rect 2844 176 2852 184
rect 3020 176 3028 184
rect 3244 176 3252 184
rect 3756 176 3764 184
rect 3948 176 3956 184
rect 4028 176 4036 184
rect 4156 176 4164 184
rect 4364 176 4372 184
rect 4716 176 4724 184
rect 4812 176 4820 184
rect 4844 176 4852 184
rect 5116 176 5124 184
rect 5164 176 5172 184
rect 5212 176 5220 184
rect 5468 176 5476 184
rect 5660 176 5668 184
rect 5916 176 5924 184
rect 6284 176 6292 184
rect 6476 176 6484 184
rect 6492 176 6500 184
rect 6684 176 6692 184
rect 7052 176 7060 184
rect 12 156 20 164
rect 44 156 52 164
rect 156 156 164 164
rect 348 156 356 164
rect 412 156 420 164
rect 572 156 580 164
rect 684 156 692 164
rect 748 156 756 164
rect 796 156 804 164
rect 876 156 884 164
rect 1004 156 1012 164
rect 1308 156 1316 164
rect 1548 156 1556 164
rect 1628 156 1636 164
rect 1708 156 1716 164
rect 1740 156 1748 164
rect 1756 156 1764 164
rect 1804 156 1812 164
rect 1820 156 1828 164
rect 1964 156 1972 164
rect 2076 156 2084 164
rect 2188 156 2196 164
rect 2252 156 2260 164
rect 2412 156 2420 164
rect 2668 156 2676 164
rect 2684 156 2692 164
rect 2716 156 2724 164
rect 2732 156 2740 164
rect 2764 156 2772 164
rect 2972 156 2980 164
rect 3036 156 3044 164
rect 3484 156 3492 164
rect 3660 156 3668 164
rect 3996 156 4004 164
rect 4012 156 4020 164
rect 4172 156 4180 164
rect 4380 156 4388 164
rect 4396 156 4404 164
rect 4764 156 4772 164
rect 5052 156 5060 164
rect 5276 156 5284 164
rect 5676 156 5684 164
rect 6092 156 6100 164
rect 92 136 100 144
rect 252 132 260 140
rect 284 136 292 144
rect 316 136 324 144
rect 508 136 516 144
rect 604 136 612 144
rect 860 136 868 144
rect 908 136 916 144
rect 940 136 948 144
rect 1020 136 1028 144
rect 1132 136 1140 144
rect 1228 136 1236 144
rect 1244 136 1252 144
rect 1436 136 1444 144
rect 1532 136 1540 144
rect 1596 136 1604 144
rect 1884 136 1892 144
rect 1900 136 1908 144
rect 1996 136 2004 144
rect 2028 136 2036 144
rect 2156 136 2164 144
rect 2284 136 2292 144
rect 2316 136 2324 144
rect 2396 136 2404 144
rect 2476 136 2484 144
rect 2588 136 2596 144
rect 2620 136 2628 144
rect 2652 136 2660 144
rect 2780 136 2788 144
rect 76 116 84 124
rect 124 116 132 124
rect 444 116 452 124
rect 492 116 500 124
rect 524 116 532 124
rect 732 116 740 124
rect 860 116 868 124
rect 1116 116 1124 124
rect 1628 116 1636 124
rect 1676 116 1684 124
rect 1740 116 1748 124
rect 1788 116 1796 124
rect 1852 116 1860 124
rect 1868 116 1876 124
rect 1932 116 1940 124
rect 1980 116 1988 124
rect 2108 116 2116 124
rect 2140 116 2148 124
rect 2236 116 2244 124
rect 2348 116 2356 124
rect 2524 116 2532 124
rect 2860 136 2868 144
rect 3004 136 3012 144
rect 3724 136 3732 144
rect 3836 136 3844 144
rect 3964 136 3972 144
rect 4044 136 4052 144
rect 4076 136 4084 144
rect 4268 136 4276 144
rect 4412 136 4420 144
rect 4556 136 4564 144
rect 4572 136 4580 144
rect 4636 136 4644 144
rect 4684 136 4692 144
rect 4700 136 4708 144
rect 4748 136 4756 144
rect 4796 136 4804 144
rect 5004 136 5012 144
rect 5036 136 5044 144
rect 5068 136 5076 144
rect 5116 136 5124 144
rect 5180 136 5188 144
rect 5244 136 5252 144
rect 5276 136 5284 144
rect 5708 136 5716 144
rect 6012 136 6020 144
rect 6092 136 6100 144
rect 6652 136 6660 144
rect 6844 136 6852 144
rect 6892 136 6900 144
rect 7196 136 7204 144
rect 7340 136 7348 144
rect 2604 116 2612 124
rect 2636 116 2644 124
rect 2684 116 2692 124
rect 2764 116 2772 124
rect 2796 116 2804 124
rect 2812 116 2820 124
rect 2908 116 2916 124
rect 3052 116 3060 124
rect 3132 116 3140 124
rect 3148 116 3156 124
rect 3228 116 3236 124
rect 3372 118 3380 126
rect 3500 116 3508 124
rect 3628 116 3636 124
rect 3676 116 3684 124
rect 3852 116 3860 124
rect 4076 116 4084 124
rect 4124 116 4132 124
rect 4252 116 4260 124
rect 4492 116 4500 124
rect 4508 116 4516 124
rect 4604 116 4612 124
rect 4652 116 4660 124
rect 4972 118 4980 126
rect 5228 116 5236 124
rect 5276 116 5284 124
rect 5340 118 5348 126
rect 5404 116 5412 124
rect 5548 116 5556 124
rect 5580 116 5588 124
rect 5692 116 5700 124
rect 5724 116 5732 124
rect 5788 118 5796 126
rect 5852 116 5860 124
rect 5996 116 6004 124
rect 6060 116 6068 124
rect 6156 118 6164 126
rect 6220 116 6228 124
rect 6396 116 6404 124
rect 6412 116 6420 124
rect 6620 118 6628 126
rect 6812 118 6820 126
rect 6940 116 6948 124
rect 7068 116 7076 124
rect 7212 116 7220 124
rect 28 96 36 104
rect 204 96 212 104
rect 284 96 292 104
rect 316 96 324 104
rect 364 96 372 104
rect 460 96 468 104
rect 604 96 612 104
rect 636 96 644 104
rect 1276 96 1284 104
rect 1692 96 1700 104
rect 2316 96 2324 104
rect 3756 96 3764 104
rect 3996 96 4004 104
rect 4108 96 4116 104
rect 4588 96 4596 104
rect 4732 96 4740 104
rect 4796 96 4804 104
rect 4828 96 4836 104
rect 5068 96 5076 104
rect 5116 96 5124 104
rect 5164 96 5172 104
rect 5212 96 5220 104
rect 6044 96 6052 104
rect 396 76 404 84
rect 444 76 452 84
rect 1468 76 1476 84
rect 1660 76 1668 84
rect 2284 76 2292 84
rect 3612 76 3620 84
rect 556 36 564 44
rect 700 36 708 44
rect 2204 36 2212 44
rect 2492 36 2500 44
rect 2540 36 2548 44
rect 3084 36 3092 44
rect 3100 36 3108 44
rect 3180 36 3188 44
rect 3196 36 3204 44
rect 3708 36 3716 44
rect 1411 6 1419 14
rect 1421 6 1429 14
rect 1431 6 1439 14
rect 1441 6 1449 14
rect 1451 6 1459 14
rect 1461 6 1469 14
rect 4419 6 4427 14
rect 4429 6 4437 14
rect 4439 6 4447 14
rect 4449 6 4457 14
rect 4459 6 4467 14
rect 4469 6 4477 14
<< metal2 >>
rect 589 5457 611 5463
rect 1245 5457 1267 5463
rect 1533 5457 1555 5463
rect 2557 5457 2579 5463
rect 605 5384 611 5457
rect 109 5304 115 5316
rect 13 5284 19 5296
rect 157 5244 163 5316
rect 253 5264 259 5356
rect 317 5344 323 5356
rect 397 5344 403 5356
rect 365 5323 371 5336
rect 461 5324 467 5376
rect 493 5344 499 5356
rect 365 5317 380 5323
rect 525 5323 531 5356
rect 541 5344 547 5356
rect 573 5324 579 5336
rect 525 5317 547 5323
rect 61 5104 67 5236
rect 141 5144 147 5236
rect 157 5123 163 5236
rect 141 5117 163 5123
rect 141 5104 147 5117
rect 157 5104 163 5117
rect 237 5104 243 5236
rect 13 5084 19 5096
rect 109 5084 115 5096
rect 76 5064 84 5070
rect 125 5064 131 5076
rect 237 5064 243 5076
rect 253 5064 259 5256
rect 301 5124 307 5236
rect 317 5224 323 5316
rect 301 5064 307 5076
rect 61 4984 67 5036
rect 77 4984 83 5036
rect 13 4744 19 4936
rect 45 4704 51 4736
rect 109 4664 115 4916
rect 125 4744 131 4936
rect 141 4924 147 4936
rect 173 4924 179 5036
rect 205 4984 211 5036
rect 253 4964 259 4976
rect 317 4963 323 5216
rect 349 5044 355 5136
rect 381 5104 387 5116
rect 397 5104 403 5236
rect 413 5104 419 5136
rect 461 5104 467 5236
rect 525 5104 531 5116
rect 397 5084 403 5096
rect 493 5064 499 5096
rect 541 5084 547 5317
rect 653 5284 659 5316
rect 669 5264 675 5336
rect 749 5324 755 5336
rect 701 5304 707 5316
rect 813 5244 819 5356
rect 845 5264 851 5316
rect 893 5264 899 5356
rect 957 5344 963 5356
rect 909 5324 915 5336
rect 973 5264 979 5316
rect 557 5124 563 5236
rect 301 4957 323 4963
rect 141 4664 147 4736
rect 157 4724 163 4916
rect 173 4904 179 4916
rect 189 4724 195 4836
rect 205 4664 211 4736
rect 13 4564 19 4636
rect 125 4564 131 4636
rect 13 4524 19 4556
rect 125 4524 131 4556
rect 189 4544 195 4636
rect 221 4624 227 4916
rect 237 4764 243 4836
rect 253 4704 259 4936
rect 301 4924 307 4957
rect 317 4904 323 4936
rect 365 4924 371 5036
rect 493 5024 499 5036
rect 397 4924 403 4976
rect 509 4944 515 5076
rect 493 4924 499 4936
rect 525 4923 531 4996
rect 589 4964 595 5096
rect 605 5084 611 5116
rect 685 5104 691 5116
rect 637 5084 643 5096
rect 605 5004 611 5036
rect 685 4984 691 5096
rect 813 5084 819 5236
rect 861 5184 867 5236
rect 941 5104 947 5236
rect 861 5097 876 5103
rect 829 5084 835 5096
rect 733 5064 739 5076
rect 861 5044 867 5097
rect 893 5044 899 5056
rect 605 4944 611 4956
rect 573 4924 579 4936
rect 621 4924 627 4936
rect 781 4924 787 5036
rect 813 4964 819 5036
rect 509 4917 531 4923
rect 253 4664 259 4696
rect 333 4584 339 4656
rect 349 4644 355 4916
rect 509 4904 515 4917
rect 733 4844 739 4916
rect 765 4904 771 4916
rect 365 4744 371 4836
rect 429 4804 435 4836
rect 365 4684 371 4736
rect 381 4663 387 4696
rect 372 4657 387 4663
rect 317 4564 323 4576
rect 333 4543 339 4576
rect 397 4564 403 4616
rect 477 4584 483 4716
rect 509 4684 515 4756
rect 557 4704 563 4756
rect 573 4684 579 4696
rect 589 4664 595 4756
rect 733 4744 739 4836
rect 669 4664 675 4676
rect 733 4664 739 4736
rect 797 4724 803 4836
rect 813 4684 819 4936
rect 861 4924 867 5036
rect 893 4963 899 5036
rect 884 4957 899 4963
rect 893 4724 899 4836
rect 893 4704 899 4716
rect 861 4697 876 4703
rect 804 4677 812 4683
rect 493 4624 499 4636
rect 445 4564 451 4576
rect 397 4544 403 4556
rect 333 4537 348 4543
rect 301 4524 307 4536
rect 429 4524 435 4556
rect 493 4524 499 4556
rect 125 4344 131 4436
rect 157 4384 163 4496
rect 125 4317 140 4323
rect 45 4264 51 4280
rect 125 4264 131 4317
rect 205 4323 211 4516
rect 205 4317 220 4323
rect 237 4264 243 4336
rect 269 4284 275 4336
rect 13 3964 19 4236
rect 61 4104 67 4196
rect 109 4144 115 4176
rect 45 3944 51 4036
rect 93 3984 99 4076
rect 13 3884 19 3936
rect 125 3924 131 4036
rect 61 3904 67 3916
rect 157 3904 163 4156
rect 205 4044 211 4116
rect 221 4104 227 4116
rect 237 4104 243 4196
rect 253 4104 259 4236
rect 285 4124 291 4296
rect 237 3984 243 4036
rect 253 3924 259 4096
rect 285 3904 291 4036
rect 29 3484 35 3636
rect 13 3404 19 3456
rect 13 3364 19 3396
rect 45 3364 51 3836
rect 93 3784 99 3896
rect 125 3884 131 3896
rect 237 3884 243 3896
rect 285 3884 291 3896
rect 253 3877 268 3883
rect 237 3864 243 3876
rect 189 3784 195 3816
rect 221 3764 227 3836
rect 253 3784 259 3877
rect 301 3864 307 3876
rect 253 3764 259 3776
rect 269 3764 275 3856
rect 317 3824 323 3896
rect 333 3844 339 4436
rect 509 4404 515 4636
rect 525 4564 531 4636
rect 621 4564 627 4656
rect 589 4524 595 4556
rect 573 4484 579 4496
rect 349 4264 355 4336
rect 365 4304 371 4316
rect 509 4284 515 4396
rect 557 4324 563 4436
rect 605 4364 611 4436
rect 621 4344 627 4516
rect 637 4504 643 4596
rect 653 4384 659 4636
rect 717 4624 723 4656
rect 701 4564 707 4596
rect 717 4584 723 4616
rect 749 4523 755 4636
rect 765 4604 771 4636
rect 797 4563 803 4676
rect 813 4624 819 4656
rect 797 4557 812 4563
rect 765 4544 771 4556
rect 845 4544 851 4576
rect 845 4524 851 4536
rect 749 4517 764 4523
rect 669 4344 675 4516
rect 669 4324 675 4336
rect 749 4324 755 4436
rect 749 4304 755 4316
rect 861 4304 867 4697
rect 893 4564 899 4676
rect 909 4664 915 4956
rect 925 4904 931 5096
rect 957 5083 963 5096
rect 948 5077 963 5083
rect 973 4984 979 5136
rect 989 5124 995 5316
rect 1005 5304 1011 5316
rect 1021 5244 1027 5336
rect 1037 5324 1043 5396
rect 1101 5384 1107 5396
rect 1261 5384 1267 5457
rect 1549 5384 1555 5457
rect 1085 5344 1091 5356
rect 1325 5344 1331 5376
rect 1485 5364 1491 5376
rect 1069 5324 1075 5336
rect 1165 5224 1171 5316
rect 1181 5304 1187 5316
rect 1053 5104 1059 5116
rect 1021 5064 1027 5096
rect 1117 5084 1123 5176
rect 1165 5164 1171 5216
rect 1149 5124 1155 5156
rect 1229 5144 1235 5316
rect 1357 5264 1363 5336
rect 1325 5184 1331 5236
rect 1165 5124 1171 5136
rect 1197 5117 1235 5123
rect 1197 5104 1203 5117
rect 1229 5104 1235 5117
rect 1165 5083 1171 5096
rect 1357 5084 1363 5256
rect 1405 5244 1411 5356
rect 1565 5344 1571 5356
rect 1373 5104 1379 5236
rect 1434 5214 1446 5216
rect 1419 5206 1421 5214
rect 1429 5206 1431 5214
rect 1439 5206 1441 5214
rect 1449 5206 1451 5214
rect 1459 5206 1461 5214
rect 1434 5204 1446 5206
rect 1485 5144 1491 5276
rect 1156 5077 1171 5083
rect 989 4964 995 5036
rect 1005 4984 1011 5016
rect 1037 4924 1043 5076
rect 1069 5024 1075 5056
rect 1133 4964 1139 5076
rect 1245 5004 1251 5036
rect 1261 4964 1267 5056
rect 1204 4957 1219 4963
rect 973 4904 979 4916
rect 1053 4764 1059 4936
rect 1149 4924 1155 4956
rect 1213 4943 1219 4957
rect 1213 4937 1228 4943
rect 1101 4784 1107 4916
rect 1245 4904 1251 4916
rect 1261 4884 1267 4956
rect 1293 4944 1299 4976
rect 1277 4924 1283 4936
rect 1309 4904 1315 4976
rect 1325 4864 1331 4876
rect 989 4704 995 4736
rect 1053 4724 1059 4736
rect 1005 4704 1011 4716
rect 957 4664 963 4676
rect 941 4644 947 4656
rect 1005 4644 1011 4676
rect 925 4583 931 4636
rect 925 4577 947 4583
rect 941 4524 947 4577
rect 973 4564 979 4636
rect 1053 4624 1059 4636
rect 1085 4584 1091 4716
rect 1101 4704 1107 4756
rect 1181 4664 1187 4676
rect 1021 4544 1027 4576
rect 1037 4523 1043 4556
rect 1085 4544 1091 4576
rect 1117 4564 1123 4656
rect 1165 4544 1171 4596
rect 1197 4584 1203 4836
rect 1357 4744 1363 4996
rect 1373 4884 1379 4896
rect 1405 4864 1411 5036
rect 1437 4964 1443 5136
rect 1517 5104 1523 5316
rect 1613 5264 1619 5356
rect 1645 5344 1651 5356
rect 1693 5324 1699 5336
rect 1661 5304 1667 5316
rect 1620 5257 1635 5263
rect 1597 5104 1603 5136
rect 1485 4984 1491 5096
rect 1501 4964 1507 5076
rect 1629 5064 1635 5257
rect 1709 5244 1715 5336
rect 1757 5244 1763 5336
rect 1917 5324 1923 5376
rect 1965 5344 1971 5356
rect 1972 5337 1987 5343
rect 1933 5324 1939 5336
rect 1789 5304 1795 5316
rect 1805 5284 1811 5296
rect 1821 5204 1827 5236
rect 1805 5103 1811 5176
rect 1869 5164 1875 5316
rect 1981 5304 1987 5337
rect 1837 5104 1843 5136
rect 1805 5097 1827 5103
rect 1517 4984 1523 5036
rect 1421 4864 1427 4956
rect 1437 4924 1443 4956
rect 1517 4944 1523 4956
rect 1597 4943 1603 5056
rect 1645 5044 1651 5096
rect 1613 4964 1619 5036
rect 1661 4964 1667 5096
rect 1789 5084 1795 5096
rect 1677 4964 1683 5056
rect 1597 4937 1612 4943
rect 1434 4814 1446 4816
rect 1419 4806 1421 4814
rect 1429 4806 1431 4814
rect 1439 4806 1441 4814
rect 1449 4806 1451 4814
rect 1459 4806 1461 4814
rect 1434 4804 1446 4806
rect 1469 4724 1475 4776
rect 1357 4704 1363 4716
rect 1277 4683 1283 4696
rect 1293 4684 1299 4696
rect 1252 4677 1283 4683
rect 1341 4664 1347 4676
rect 1213 4604 1219 4636
rect 1293 4543 1299 4636
rect 1284 4537 1299 4543
rect 1037 4517 1052 4523
rect 1053 4504 1059 4516
rect 365 4164 371 4236
rect 381 4164 387 4256
rect 413 4244 419 4276
rect 509 4264 515 4276
rect 605 4264 611 4276
rect 413 4124 419 4236
rect 461 4204 467 4236
rect 541 4164 547 4236
rect 701 4204 707 4296
rect 877 4284 883 4436
rect 893 4324 899 4436
rect 925 4324 931 4376
rect 989 4344 995 4436
rect 973 4304 979 4316
rect 749 4264 755 4276
rect 861 4244 867 4276
rect 893 4244 899 4296
rect 925 4284 931 4296
rect 989 4284 995 4336
rect 1069 4324 1075 4436
rect 1149 4344 1155 4396
rect 1149 4324 1155 4336
rect 1053 4304 1059 4316
rect 397 3944 403 4036
rect 429 4024 435 4136
rect 477 3904 483 3916
rect 461 3864 467 3876
rect 349 3756 355 3836
rect 413 3744 419 3836
rect 477 3784 483 3896
rect 429 3744 435 3776
rect 509 3764 515 3796
rect 525 3764 531 3876
rect 557 3764 563 4076
rect 605 4044 611 4136
rect 621 3944 627 4156
rect 637 4024 643 4136
rect 781 4124 787 4216
rect 829 4164 835 4236
rect 621 3884 627 3936
rect 637 3917 652 3923
rect 573 3864 579 3876
rect 637 3864 643 3917
rect 685 3884 691 3936
rect 733 3824 739 3856
rect 621 3764 627 3796
rect 477 3744 483 3756
rect 717 3744 723 3756
rect 109 3724 115 3736
rect 141 3703 147 3736
rect 237 3724 243 3736
rect 557 3724 563 3736
rect 605 3724 611 3736
rect 141 3697 163 3703
rect 61 3504 67 3576
rect 77 3364 83 3476
rect 125 3424 131 3456
rect 13 3024 19 3056
rect 13 2964 19 3016
rect 61 2924 67 3096
rect 77 3064 83 3316
rect 109 3304 115 3316
rect 157 3263 163 3697
rect 173 3504 179 3576
rect 173 3464 179 3496
rect 205 3483 211 3636
rect 285 3504 291 3576
rect 317 3504 323 3676
rect 205 3477 220 3483
rect 173 3424 179 3436
rect 173 3284 179 3316
rect 157 3257 179 3263
rect 109 3144 115 3236
rect 93 2924 99 2936
rect 61 2704 67 2916
rect 109 2904 115 3116
rect 141 3044 147 3076
rect 157 3024 163 3056
rect 141 2944 147 2976
rect 109 2724 115 2896
rect 13 2604 19 2656
rect 13 2564 19 2596
rect 61 2524 67 2696
rect 93 2684 99 2696
rect 109 2504 115 2716
rect 141 2644 147 2676
rect 157 2604 163 2656
rect 141 2544 147 2576
rect 157 2564 163 2596
rect 173 2543 179 3257
rect 205 3104 211 3456
rect 237 3424 243 3456
rect 253 3124 259 3496
rect 285 3364 291 3436
rect 301 3364 307 3476
rect 333 3344 339 3536
rect 349 3463 355 3636
rect 557 3584 563 3716
rect 589 3704 595 3716
rect 413 3504 419 3536
rect 461 3504 467 3536
rect 509 3524 515 3536
rect 349 3457 364 3463
rect 541 3444 547 3476
rect 621 3464 627 3636
rect 669 3503 675 3636
rect 660 3497 675 3503
rect 685 3464 691 3596
rect 701 3504 707 3516
rect 717 3483 723 3716
rect 733 3604 739 3636
rect 749 3583 755 4036
rect 765 3884 771 3896
rect 765 3744 771 3816
rect 797 3803 803 4116
rect 861 4004 867 4156
rect 909 4123 915 4276
rect 925 4197 988 4203
rect 925 4164 931 4197
rect 1005 4184 1011 4276
rect 1037 4184 1043 4236
rect 1053 4184 1059 4216
rect 1021 4164 1027 4176
rect 1085 4144 1091 4296
rect 1133 4244 1139 4256
rect 1117 4164 1123 4196
rect 957 4124 963 4136
rect 900 4117 915 4123
rect 909 4064 915 4117
rect 1044 4117 1068 4123
rect 1005 4084 1011 4096
rect 1085 4084 1091 4116
rect 1133 4084 1139 4236
rect 861 3884 867 3936
rect 877 3904 883 4036
rect 813 3824 819 3876
rect 845 3864 851 3876
rect 877 3864 883 3896
rect 797 3797 819 3803
rect 701 3477 723 3483
rect 733 3577 755 3583
rect 733 3483 739 3577
rect 797 3564 803 3636
rect 813 3624 819 3797
rect 829 3724 835 3816
rect 845 3764 851 3856
rect 845 3744 851 3756
rect 861 3744 867 3836
rect 893 3744 899 3956
rect 909 3863 915 4016
rect 925 3884 931 3896
rect 1069 3884 1075 4036
rect 1101 3984 1107 3996
rect 1117 3923 1123 4076
rect 1101 3917 1123 3923
rect 1021 3864 1027 3876
rect 909 3857 931 3863
rect 909 3804 915 3836
rect 749 3524 755 3556
rect 813 3504 819 3516
rect 765 3484 771 3496
rect 733 3477 748 3483
rect 333 3324 339 3336
rect 381 3324 387 3436
rect 493 3404 499 3436
rect 413 3164 419 3316
rect 429 3284 435 3336
rect 477 3284 483 3316
rect 493 3284 499 3376
rect 509 3304 515 3436
rect 557 3324 563 3356
rect 253 3104 259 3116
rect 269 3084 275 3096
rect 253 3064 259 3076
rect 205 2964 211 2996
rect 269 2944 275 2956
rect 285 2944 291 3036
rect 317 3024 323 3056
rect 205 2704 211 2836
rect 237 2704 243 2856
rect 253 2844 259 2916
rect 285 2864 291 2916
rect 205 2544 211 2696
rect 157 2537 179 2543
rect 61 2303 67 2436
rect 109 2304 115 2316
rect 52 2297 67 2303
rect 29 2124 35 2236
rect 77 2224 83 2256
rect 77 2124 83 2156
rect 93 2144 99 2276
rect 125 2264 131 2276
rect 141 2144 147 2176
rect 13 1984 19 2096
rect 45 2084 51 2116
rect 141 2064 147 2116
rect 61 1924 67 2036
rect 13 1884 19 1896
rect 141 1884 147 1896
rect 109 1864 115 1876
rect 45 1803 51 1856
rect 61 1824 67 1856
rect 45 1797 67 1803
rect 13 1764 19 1796
rect 61 1784 67 1797
rect 125 1764 131 1796
rect 141 1743 147 1856
rect 157 1844 163 2537
rect 189 2224 195 2256
rect 205 2224 211 2256
rect 173 2104 179 2136
rect 189 1984 195 2116
rect 205 2104 211 2136
rect 221 2124 227 2516
rect 237 2324 243 2536
rect 237 2304 243 2316
rect 253 2164 259 2316
rect 285 2304 291 2856
rect 333 2684 339 3116
rect 349 2904 355 3136
rect 365 2924 371 2936
rect 397 2844 403 3096
rect 477 3064 483 3236
rect 509 3064 515 3096
rect 413 2964 419 3056
rect 445 3024 451 3056
rect 461 3044 467 3056
rect 477 2943 483 3036
rect 461 2937 483 2943
rect 349 2704 355 2816
rect 349 2644 355 2676
rect 365 2624 371 2836
rect 413 2723 419 2936
rect 445 2883 451 2916
rect 461 2904 467 2937
rect 493 2884 499 2956
rect 525 2944 531 2976
rect 445 2877 467 2883
rect 461 2784 467 2877
rect 397 2717 419 2723
rect 397 2684 403 2717
rect 461 2704 467 2756
rect 397 2564 403 2676
rect 413 2664 419 2696
rect 317 2524 323 2536
rect 381 2524 387 2536
rect 461 2524 467 2536
rect 317 2144 323 2436
rect 381 2363 387 2436
rect 365 2357 387 2363
rect 365 2324 371 2357
rect 461 2324 467 2436
rect 493 2364 499 2816
rect 509 2784 515 2836
rect 525 2824 531 2916
rect 509 2704 515 2716
rect 509 2544 515 2696
rect 525 2484 531 2736
rect 541 2723 547 3236
rect 589 3084 595 3096
rect 605 3063 611 3436
rect 621 3104 627 3316
rect 637 3304 643 3436
rect 653 3084 659 3396
rect 669 3344 675 3436
rect 701 3324 707 3477
rect 749 3464 755 3476
rect 717 3324 723 3436
rect 765 3324 771 3336
rect 781 3324 787 3396
rect 797 3364 803 3436
rect 813 3404 819 3436
rect 669 3284 675 3316
rect 740 3297 755 3303
rect 669 3084 675 3276
rect 701 3224 707 3276
rect 717 3103 723 3236
rect 708 3097 723 3103
rect 733 3084 739 3276
rect 749 3244 755 3297
rect 804 3297 819 3303
rect 765 3264 771 3276
rect 765 3064 771 3196
rect 813 3184 819 3297
rect 605 3057 620 3063
rect 637 2964 643 3036
rect 589 2924 595 2956
rect 621 2744 627 2956
rect 669 2903 675 3036
rect 717 2964 723 3036
rect 749 2924 755 3036
rect 765 2924 771 2976
rect 653 2897 675 2903
rect 653 2764 659 2897
rect 541 2717 556 2723
rect 669 2704 675 2836
rect 701 2804 707 2896
rect 717 2703 723 2856
rect 765 2724 771 2876
rect 781 2784 787 2796
rect 797 2764 803 3136
rect 813 3104 819 3156
rect 813 2924 819 2936
rect 829 2903 835 3676
rect 845 3484 851 3716
rect 877 3704 883 3716
rect 877 3504 883 3696
rect 925 3504 931 3857
rect 957 3764 963 3796
rect 941 3564 947 3756
rect 973 3744 979 3816
rect 989 3784 995 3836
rect 1037 3784 1043 3836
rect 1069 3744 1075 3856
rect 1085 3744 1091 3916
rect 1101 3784 1107 3917
rect 1117 3884 1123 3896
rect 1133 3864 1139 4036
rect 1149 4024 1155 4036
rect 1165 4004 1171 4536
rect 1181 4504 1187 4536
rect 1277 4517 1292 4523
rect 1229 4324 1235 4436
rect 1181 4264 1187 4276
rect 1181 4124 1187 4136
rect 1181 3923 1187 3936
rect 1197 3923 1203 4036
rect 1181 3917 1203 3923
rect 1181 3904 1187 3917
rect 1213 3904 1219 4276
rect 1229 4124 1235 4216
rect 1261 4164 1267 4296
rect 1277 4224 1283 4517
rect 1309 4523 1315 4616
rect 1300 4517 1315 4523
rect 1325 4364 1331 4536
rect 1341 4323 1347 4436
rect 1357 4344 1363 4696
rect 1517 4684 1523 4696
rect 1533 4684 1539 4836
rect 1581 4744 1587 4936
rect 1613 4824 1619 4936
rect 1661 4844 1667 4956
rect 1709 4944 1715 5076
rect 1805 5064 1811 5076
rect 1773 5024 1779 5036
rect 1757 4984 1763 4996
rect 1821 4984 1827 5097
rect 1853 5064 1859 5076
rect 1821 4944 1827 4976
rect 1853 4964 1859 5056
rect 1869 5024 1875 5116
rect 1885 4944 1891 5076
rect 1901 5064 1907 5096
rect 1917 5084 1923 5176
rect 1933 5124 1939 5136
rect 1908 5057 1923 5063
rect 1901 4944 1907 4956
rect 1837 4924 1843 4936
rect 1869 4924 1875 4936
rect 1917 4924 1923 5057
rect 1949 4904 1955 5036
rect 1965 4964 1971 5076
rect 1981 5064 1987 5296
rect 2013 5244 2019 5356
rect 2029 5344 2035 5376
rect 2333 5364 2339 5376
rect 2077 5324 2083 5356
rect 2109 5344 2115 5356
rect 2205 5344 2211 5356
rect 2381 5344 2387 5356
rect 2093 5324 2099 5336
rect 2205 5324 2211 5336
rect 2093 5304 2099 5316
rect 2013 5184 2019 5236
rect 2045 5084 2051 5176
rect 2061 5104 2067 5236
rect 2093 5064 2099 5256
rect 2109 5104 2115 5196
rect 2141 5123 2147 5316
rect 2157 5264 2163 5296
rect 2173 5284 2179 5316
rect 2221 5304 2227 5336
rect 2317 5324 2323 5336
rect 2525 5324 2531 5336
rect 2269 5204 2275 5316
rect 2269 5184 2275 5196
rect 2365 5184 2371 5236
rect 2189 5137 2204 5143
rect 2141 5117 2156 5123
rect 2157 5084 2163 5096
rect 1997 4964 2003 5016
rect 1965 4924 1971 4956
rect 1981 4864 1987 4916
rect 2029 4903 2035 5036
rect 2045 4924 2051 5016
rect 2077 4984 2083 5036
rect 2029 4897 2044 4903
rect 2029 4864 2035 4876
rect 1837 4704 1843 4836
rect 1405 4544 1411 4556
rect 1332 4317 1347 4323
rect 1293 4284 1299 4316
rect 1325 4284 1331 4316
rect 1373 4304 1379 4476
rect 1389 4384 1395 4536
rect 1434 4414 1446 4416
rect 1419 4406 1421 4414
rect 1429 4406 1431 4414
rect 1439 4406 1441 4414
rect 1449 4406 1451 4414
rect 1459 4406 1461 4414
rect 1434 4404 1446 4406
rect 1421 4304 1427 4376
rect 1485 4363 1491 4636
rect 1501 4384 1507 4536
rect 1549 4523 1555 4636
rect 1565 4604 1571 4656
rect 1597 4564 1603 4636
rect 1613 4544 1619 4556
rect 1629 4544 1635 4676
rect 1725 4644 1731 4676
rect 1661 4524 1667 4636
rect 1741 4564 1747 4696
rect 1789 4684 1795 4696
rect 1837 4684 1843 4696
rect 1933 4684 1939 4816
rect 1933 4664 1939 4676
rect 1757 4584 1763 4596
rect 1853 4584 1859 4636
rect 1917 4584 1923 4596
rect 1933 4563 1939 4656
rect 1949 4624 1955 4696
rect 1965 4584 1971 4676
rect 1981 4584 1987 4836
rect 1997 4684 2003 4696
rect 1917 4557 1939 4563
rect 1709 4524 1715 4556
rect 1549 4517 1571 4523
rect 1485 4357 1507 4363
rect 1437 4284 1443 4356
rect 1309 4144 1315 4156
rect 1277 4124 1283 4136
rect 1325 4104 1331 4236
rect 1373 4164 1379 4276
rect 1389 4123 1395 4236
rect 1405 4164 1411 4216
rect 1437 4144 1443 4196
rect 1380 4117 1395 4123
rect 1277 3904 1283 4056
rect 1373 3944 1379 4036
rect 1485 4024 1491 4336
rect 1501 4284 1507 4357
rect 1565 4324 1571 4517
rect 1709 4384 1715 4516
rect 1757 4463 1763 4496
rect 1757 4457 1779 4463
rect 1613 4304 1619 4376
rect 1629 4284 1635 4336
rect 1501 4164 1507 4276
rect 1581 4144 1587 4236
rect 1629 4184 1635 4276
rect 1661 4264 1667 4356
rect 1709 4244 1715 4296
rect 1725 4284 1731 4316
rect 1741 4284 1747 4296
rect 1741 4264 1747 4276
rect 1645 4224 1651 4236
rect 1709 4144 1715 4156
rect 1773 4144 1779 4457
rect 1789 4304 1795 4336
rect 1821 4284 1827 4516
rect 1869 4364 1875 4556
rect 1901 4523 1907 4536
rect 1917 4523 1923 4557
rect 2013 4544 2019 4736
rect 2045 4563 2051 4836
rect 2077 4824 2083 4956
rect 2109 4944 2115 5056
rect 2157 4944 2163 5036
rect 2173 5004 2179 5116
rect 2189 4944 2195 5137
rect 2205 5104 2211 5136
rect 2285 5104 2291 5116
rect 2429 5104 2435 5116
rect 2477 5104 2483 5136
rect 2228 5077 2243 5083
rect 2221 4964 2227 4996
rect 2237 4984 2243 5077
rect 2237 4924 2243 4976
rect 2269 4924 2275 5036
rect 2317 4964 2323 5036
rect 2333 5004 2339 5056
rect 2365 4964 2371 5056
rect 2381 4964 2387 5076
rect 2413 4964 2419 5076
rect 2365 4924 2371 4956
rect 2381 4944 2387 4956
rect 2461 4944 2467 4956
rect 2477 4944 2483 5056
rect 2493 4984 2499 5236
rect 2525 5184 2531 5296
rect 2541 5184 2547 5316
rect 2557 5304 2563 5416
rect 2573 5384 2579 5457
rect 2589 5424 2595 5463
rect 2797 5457 2819 5463
rect 2845 5457 2867 5463
rect 2813 5384 2819 5457
rect 2861 5384 2867 5457
rect 3005 5457 3027 5463
rect 2938 5414 2950 5416
rect 2923 5406 2925 5414
rect 2933 5406 2935 5414
rect 2943 5406 2945 5414
rect 2953 5406 2955 5414
rect 2963 5406 2965 5414
rect 2938 5404 2950 5406
rect 2589 5344 2595 5376
rect 2685 5304 2691 5356
rect 2589 5024 2595 5036
rect 2541 4984 2547 4996
rect 2605 4964 2611 5076
rect 2637 4984 2643 4996
rect 2509 4924 2515 4936
rect 2173 4903 2179 4916
rect 2164 4897 2179 4903
rect 2461 4903 2467 4916
rect 2461 4897 2476 4903
rect 2509 4844 2515 4916
rect 2205 4804 2211 4836
rect 2301 4784 2307 4836
rect 2061 4704 2067 4736
rect 2109 4697 2124 4703
rect 2077 4644 2083 4676
rect 2061 4564 2067 4636
rect 2109 4584 2115 4697
rect 2173 4684 2179 4716
rect 2205 4644 2211 4696
rect 2036 4557 2051 4563
rect 2077 4543 2083 4556
rect 2141 4544 2147 4556
rect 2068 4537 2083 4543
rect 1901 4517 1923 4523
rect 1917 4444 1923 4517
rect 1933 4504 1939 4536
rect 2157 4524 2163 4576
rect 1972 4517 1987 4523
rect 1933 4284 1939 4296
rect 1869 4264 1875 4276
rect 1434 4014 1446 4016
rect 1419 4006 1421 4014
rect 1429 4006 1431 4014
rect 1439 4006 1441 4014
rect 1449 4006 1451 4014
rect 1459 4006 1461 4014
rect 1434 4004 1446 4006
rect 1389 3923 1395 3996
rect 1533 3944 1539 4136
rect 1805 4124 1811 4236
rect 1853 4104 1859 4116
rect 1389 3917 1411 3923
rect 1213 3864 1219 3896
rect 1261 3884 1267 3896
rect 1389 3884 1395 3896
rect 1405 3884 1411 3917
rect 1245 3744 1251 3836
rect 1261 3723 1267 3836
rect 1469 3804 1475 3936
rect 1565 3904 1571 4036
rect 1581 3884 1587 4076
rect 1661 3943 1667 4096
rect 1885 3984 1891 4276
rect 1917 4264 1923 4276
rect 1949 4184 1955 4476
rect 1965 4204 1971 4416
rect 1981 4384 1987 4517
rect 2205 4504 2211 4556
rect 2221 4524 2227 4576
rect 1981 4304 1987 4356
rect 1949 4143 1955 4176
rect 1933 4137 1955 4143
rect 1933 4124 1939 4137
rect 1965 4123 1971 4196
rect 1997 4124 2003 4456
rect 2029 4384 2035 4436
rect 2045 4364 2051 4496
rect 2237 4484 2243 4576
rect 2253 4544 2259 4656
rect 2317 4584 2323 4696
rect 2333 4684 2339 4836
rect 2429 4724 2435 4796
rect 2365 4664 2371 4716
rect 2381 4664 2387 4696
rect 2461 4684 2467 4836
rect 2493 4704 2499 4796
rect 2509 4683 2515 4796
rect 2541 4704 2547 4736
rect 2493 4677 2515 4683
rect 2413 4664 2419 4676
rect 2349 4544 2355 4636
rect 2061 4304 2067 4336
rect 2077 4324 2083 4396
rect 2141 4304 2147 4336
rect 2157 4304 2163 4436
rect 2221 4403 2227 4436
rect 2205 4397 2227 4403
rect 2173 4324 2179 4356
rect 2189 4304 2195 4336
rect 2205 4304 2211 4397
rect 2237 4364 2243 4476
rect 2253 4384 2259 4396
rect 2269 4324 2275 4436
rect 2285 4324 2291 4536
rect 2365 4524 2371 4636
rect 2349 4424 2355 4516
rect 2381 4424 2387 4616
rect 2429 4563 2435 4636
rect 2420 4557 2435 4563
rect 2461 4544 2467 4596
rect 2493 4524 2499 4677
rect 2445 4444 2451 4516
rect 2493 4484 2499 4516
rect 2349 4364 2355 4416
rect 2397 4384 2403 4436
rect 2333 4324 2339 4336
rect 2068 4297 2083 4303
rect 1956 4117 1971 4123
rect 1661 3937 1683 3943
rect 1677 3884 1683 3937
rect 1821 3904 1827 3916
rect 1885 3904 1891 3976
rect 1949 3924 1955 3936
rect 1981 3904 1987 4096
rect 1997 3924 2003 3936
rect 1997 3904 2003 3916
rect 2013 3904 2019 4256
rect 2077 4124 2083 4297
rect 2237 4284 2243 4296
rect 2029 3984 2035 4016
rect 1565 3864 1571 3876
rect 1245 3717 1267 3723
rect 1229 3704 1235 3716
rect 1245 3704 1251 3717
rect 1284 3717 1299 3723
rect 1277 3704 1283 3716
rect 1261 3664 1267 3696
rect 1053 3584 1059 3616
rect 1021 3524 1027 3556
rect 1117 3544 1123 3556
rect 1053 3484 1059 3496
rect 909 3464 915 3476
rect 884 3317 899 3323
rect 845 3283 851 3316
rect 845 3277 860 3283
rect 877 3184 883 3236
rect 893 3083 899 3317
rect 941 3284 947 3476
rect 957 3324 963 3456
rect 973 3444 979 3456
rect 909 3144 915 3236
rect 941 3184 947 3216
rect 973 3184 979 3336
rect 989 3304 995 3436
rect 1069 3364 1075 3476
rect 1005 3284 1011 3316
rect 1021 3304 1027 3336
rect 1101 3324 1107 3496
rect 1133 3343 1139 3636
rect 1229 3563 1235 3636
rect 1277 3564 1283 3676
rect 1293 3584 1299 3717
rect 1229 3557 1251 3563
rect 1181 3524 1187 3536
rect 1181 3503 1187 3516
rect 1181 3497 1203 3503
rect 1149 3444 1155 3476
rect 1117 3337 1139 3343
rect 1053 3304 1059 3316
rect 1021 3284 1027 3296
rect 1069 3263 1075 3316
rect 1117 3304 1123 3337
rect 1149 3284 1155 3316
rect 1165 3263 1171 3496
rect 1069 3257 1091 3263
rect 1165 3257 1187 3263
rect 1021 3184 1027 3256
rect 1037 3124 1043 3236
rect 877 3077 899 3083
rect 877 2984 883 3077
rect 909 2984 915 3096
rect 925 3064 931 3096
rect 845 2944 851 2976
rect 829 2897 851 2903
rect 797 2744 803 2756
rect 813 2724 819 2896
rect 708 2697 723 2703
rect 765 2703 771 2716
rect 765 2697 780 2703
rect 541 2524 547 2676
rect 573 2644 579 2696
rect 829 2664 835 2696
rect 589 2524 595 2536
rect 605 2444 611 2636
rect 621 2624 627 2656
rect 621 2544 627 2576
rect 701 2564 707 2636
rect 717 2524 723 2656
rect 813 2584 819 2636
rect 829 2584 835 2656
rect 845 2644 851 2897
rect 877 2684 883 2796
rect 893 2784 899 2896
rect 909 2884 915 2976
rect 941 2943 947 2976
rect 957 2964 963 2996
rect 941 2937 963 2943
rect 493 2304 499 2356
rect 653 2324 659 2436
rect 669 2304 675 2356
rect 765 2344 771 2436
rect 781 2344 787 2476
rect 333 2184 339 2296
rect 413 2264 419 2296
rect 525 2284 531 2296
rect 365 2144 371 2176
rect 205 1924 211 2076
rect 180 1897 195 1903
rect 173 1864 179 1876
rect 189 1824 195 1897
rect 237 1903 243 2036
rect 237 1897 252 1903
rect 205 1804 211 1896
rect 269 1764 275 1916
rect 285 1904 291 2096
rect 317 2084 323 2096
rect 349 2044 355 2136
rect 381 2124 387 2236
rect 461 2184 467 2256
rect 477 2244 483 2276
rect 557 2184 563 2296
rect 605 2264 611 2296
rect 621 2284 627 2296
rect 781 2284 787 2336
rect 829 2304 835 2516
rect 893 2504 899 2716
rect 909 2664 915 2716
rect 925 2684 931 2796
rect 957 2684 963 2937
rect 973 2744 979 3016
rect 989 2904 995 3096
rect 1005 3084 1011 3096
rect 1005 3064 1011 3076
rect 1021 2944 1027 3076
rect 1069 3044 1075 3076
rect 1085 3024 1091 3257
rect 1101 3084 1107 3236
rect 1149 3144 1155 3156
rect 1133 3103 1139 3116
rect 1165 3104 1171 3236
rect 1124 3097 1139 3103
rect 1085 2964 1091 2996
rect 1117 2943 1123 3016
rect 1117 2937 1132 2943
rect 989 2824 995 2896
rect 1005 2884 1011 2916
rect 1005 2857 1011 2876
rect 1021 2764 1027 2936
rect 1053 2844 1059 2916
rect 1101 2884 1107 2896
rect 1085 2784 1091 2876
rect 1101 2804 1107 2876
rect 1117 2784 1123 2937
rect 1149 2924 1155 2936
rect 973 2684 979 2716
rect 1021 2684 1027 2716
rect 845 2344 851 2476
rect 909 2344 915 2636
rect 957 2604 963 2676
rect 973 2644 979 2676
rect 1005 2664 1011 2676
rect 957 2524 963 2596
rect 989 2564 995 2596
rect 1005 2584 1011 2656
rect 1037 2524 1043 2776
rect 1069 2684 1075 2716
rect 1101 2564 1107 2596
rect 1133 2524 1139 2876
rect 1181 2704 1187 3257
rect 1197 3124 1203 3497
rect 1213 3464 1219 3496
rect 1213 3384 1219 3436
rect 1229 3384 1235 3536
rect 1213 3324 1219 3336
rect 1229 3143 1235 3356
rect 1245 3343 1251 3557
rect 1277 3484 1283 3556
rect 1293 3504 1299 3576
rect 1245 3340 1267 3343
rect 1245 3337 1260 3340
rect 1277 3244 1283 3336
rect 1293 3304 1299 3436
rect 1309 3364 1315 3636
rect 1325 3584 1331 3676
rect 1325 3284 1331 3536
rect 1341 3524 1347 3736
rect 1373 3704 1379 3716
rect 1357 3644 1363 3696
rect 1373 3564 1379 3696
rect 1501 3684 1507 3696
rect 1517 3664 1523 3716
rect 1533 3704 1539 3836
rect 1565 3684 1571 3696
rect 1581 3664 1587 3716
rect 1613 3703 1619 3836
rect 1693 3824 1699 3896
rect 1901 3884 1907 3896
rect 1837 3864 1843 3876
rect 1677 3744 1683 3776
rect 1645 3704 1651 3716
rect 1604 3697 1619 3703
rect 1661 3684 1667 3696
rect 1373 3524 1379 3536
rect 1389 3504 1395 3656
rect 1434 3614 1446 3616
rect 1419 3606 1421 3614
rect 1429 3606 1431 3614
rect 1439 3606 1441 3614
rect 1449 3606 1451 3614
rect 1459 3606 1461 3614
rect 1434 3604 1446 3606
rect 1405 3544 1411 3556
rect 1341 3484 1347 3496
rect 1357 3324 1363 3336
rect 1389 3324 1395 3476
rect 1453 3384 1459 3576
rect 1517 3524 1523 3636
rect 1581 3624 1587 3636
rect 1485 3323 1491 3356
rect 1501 3344 1507 3476
rect 1485 3317 1500 3323
rect 1229 3137 1251 3143
rect 1197 3004 1203 3076
rect 1229 2944 1235 2956
rect 1197 2924 1203 2936
rect 1197 2884 1203 2896
rect 1197 2704 1203 2876
rect 1197 2664 1203 2676
rect 1181 2644 1187 2656
rect 1149 2524 1155 2636
rect 1165 2544 1171 2556
rect 845 2284 851 2336
rect 877 2304 883 2336
rect 669 2244 675 2276
rect 404 2117 419 2123
rect 413 2104 419 2117
rect 349 1984 355 1996
rect 397 1924 403 2096
rect 445 2084 451 2136
rect 493 2084 499 2176
rect 589 2144 595 2176
rect 685 2144 691 2236
rect 829 2144 835 2236
rect 845 2184 851 2216
rect 541 2104 547 2116
rect 500 2077 515 2083
rect 189 1744 195 1756
rect 125 1737 147 1743
rect 109 1704 115 1736
rect 29 1584 35 1656
rect 61 1584 67 1696
rect 125 1584 131 1737
rect 173 1724 179 1736
rect 157 1584 163 1676
rect 221 1584 227 1716
rect 237 1684 243 1736
rect 269 1664 275 1736
rect 301 1724 307 1876
rect 333 1864 339 1916
rect 413 1903 419 1916
rect 429 1904 435 1916
rect 404 1897 419 1903
rect 365 1844 371 1876
rect 445 1824 451 1936
rect 493 1924 499 1956
rect 509 1944 515 2077
rect 525 2064 531 2096
rect 541 2084 547 2096
rect 557 1984 563 2056
rect 573 1963 579 2136
rect 861 2124 867 2236
rect 628 2117 643 2123
rect 637 2104 643 2117
rect 589 1984 595 2036
rect 653 1984 659 2116
rect 733 2064 739 2116
rect 813 2084 819 2116
rect 877 2084 883 2256
rect 909 2244 915 2296
rect 925 2104 931 2236
rect 957 2224 963 2296
rect 964 2217 979 2223
rect 941 2124 947 2136
rect 573 1957 595 1963
rect 461 1917 476 1923
rect 333 1724 339 1796
rect 381 1764 387 1796
rect 397 1784 403 1816
rect 413 1724 419 1756
rect 429 1744 435 1756
rect 308 1717 323 1723
rect 285 1703 291 1716
rect 285 1697 300 1703
rect 317 1684 323 1717
rect 429 1704 435 1716
rect 461 1664 467 1917
rect 493 1884 499 1896
rect 509 1764 515 1796
rect 541 1764 547 1856
rect 573 1784 579 1896
rect 589 1784 595 1957
rect 701 1924 707 1976
rect 685 1904 691 1916
rect 685 1884 691 1896
rect 717 1884 723 1896
rect 637 1864 643 1876
rect 573 1744 579 1756
rect 477 1724 483 1736
rect 285 1584 291 1656
rect 365 1504 371 1556
rect 61 1477 76 1483
rect 13 1384 19 1456
rect 61 1364 67 1477
rect 77 1464 83 1476
rect 93 1364 99 1480
rect 141 1444 147 1456
rect 205 1444 211 1496
rect 237 1443 243 1456
rect 317 1444 323 1496
rect 237 1437 259 1443
rect 205 1364 211 1436
rect 61 1284 67 1356
rect 77 1344 83 1356
rect 93 1284 99 1316
rect 173 1264 179 1316
rect 173 1124 179 1136
rect 189 1124 195 1236
rect 205 1184 211 1336
rect 221 1324 227 1356
rect 13 1084 19 1096
rect 61 1064 67 1076
rect 157 1044 163 1076
rect 109 984 115 1036
rect 125 984 131 1036
rect 221 1004 227 1076
rect 237 1044 243 1056
rect 253 1023 259 1437
rect 365 1384 371 1496
rect 397 1484 403 1496
rect 413 1384 419 1536
rect 557 1484 563 1716
rect 573 1504 579 1736
rect 685 1584 691 1876
rect 717 1784 723 1816
rect 733 1763 739 2036
rect 765 1924 771 2036
rect 781 1763 787 1956
rect 877 1904 883 2076
rect 973 2064 979 2217
rect 989 2184 995 2476
rect 1005 2344 1011 2376
rect 1037 2364 1043 2516
rect 1197 2504 1203 2656
rect 1021 2304 1027 2316
rect 1005 2124 1011 2136
rect 909 1884 915 2036
rect 941 1984 947 2056
rect 868 1877 883 1883
rect 845 1843 851 1876
rect 861 1864 867 1876
rect 845 1837 867 1843
rect 717 1757 739 1763
rect 765 1757 787 1763
rect 701 1584 707 1736
rect 685 1544 691 1576
rect 461 1444 467 1456
rect 493 1364 499 1456
rect 509 1364 515 1436
rect 269 1184 275 1356
rect 509 1344 515 1356
rect 541 1344 547 1476
rect 557 1464 563 1476
rect 365 1324 371 1336
rect 461 1324 467 1336
rect 292 1317 348 1323
rect 365 1284 371 1316
rect 541 1304 547 1336
rect 557 1324 563 1396
rect 605 1324 611 1396
rect 653 1384 659 1436
rect 669 1404 675 1476
rect 717 1384 723 1757
rect 765 1744 771 1757
rect 861 1744 867 1837
rect 877 1764 883 1877
rect 925 1864 931 1916
rect 941 1904 947 1936
rect 957 1924 963 1936
rect 973 1904 979 2056
rect 1005 1924 1011 2036
rect 941 1784 947 1896
rect 973 1784 979 1856
rect 989 1844 995 1916
rect 1037 1864 1043 2316
rect 1069 2203 1075 2436
rect 1085 2304 1091 2376
rect 1165 2304 1171 2316
rect 1181 2284 1187 2416
rect 1213 2384 1219 2936
rect 1245 2863 1251 3137
rect 1261 2984 1267 3076
rect 1261 2924 1267 2956
rect 1277 2924 1283 3056
rect 1325 2984 1331 3116
rect 1341 3104 1347 3236
rect 1357 3124 1363 3296
rect 1373 3184 1379 3196
rect 1389 3184 1395 3316
rect 1517 3224 1523 3336
rect 1434 3214 1446 3216
rect 1419 3206 1421 3214
rect 1429 3206 1431 3214
rect 1439 3206 1441 3214
rect 1449 3206 1451 3214
rect 1459 3206 1461 3214
rect 1434 3204 1446 3206
rect 1533 3204 1539 3336
rect 1549 3324 1555 3516
rect 1597 3504 1603 3636
rect 1629 3584 1635 3676
rect 1613 3503 1619 3516
rect 1613 3497 1628 3503
rect 1597 3364 1603 3436
rect 1645 3343 1651 3636
rect 1677 3484 1683 3596
rect 1661 3444 1667 3476
rect 1693 3463 1699 3716
rect 1709 3484 1715 3516
rect 1725 3504 1731 3716
rect 1741 3504 1747 3616
rect 1693 3457 1715 3463
rect 1693 3403 1699 3436
rect 1709 3404 1715 3457
rect 1629 3337 1651 3343
rect 1677 3397 1699 3403
rect 1629 3324 1635 3337
rect 1677 3324 1683 3397
rect 1693 3344 1699 3376
rect 1709 3364 1715 3376
rect 1645 3317 1660 3323
rect 1645 3304 1651 3317
rect 1613 3264 1619 3276
rect 1581 3184 1587 3236
rect 1645 3184 1651 3216
rect 1725 3204 1731 3476
rect 1757 3464 1763 3836
rect 1773 3764 1779 3796
rect 1949 3764 1955 3796
rect 1997 3764 2003 3796
rect 1837 3704 1843 3756
rect 2013 3744 2019 3896
rect 2045 3824 2051 4036
rect 2061 3944 2067 4056
rect 2061 3904 2067 3936
rect 1917 3724 1923 3736
rect 1805 3584 1811 3676
rect 1821 3504 1827 3636
rect 1821 3384 1827 3436
rect 1773 3224 1779 3276
rect 1805 3264 1811 3296
rect 1709 3184 1715 3196
rect 1357 3083 1363 3116
rect 1421 3084 1427 3096
rect 1341 3077 1363 3083
rect 1309 2944 1315 2976
rect 1277 2884 1283 2916
rect 1245 2857 1267 2863
rect 1245 2724 1251 2796
rect 1229 2564 1235 2596
rect 1245 2564 1251 2616
rect 1101 2244 1107 2256
rect 1069 2197 1091 2203
rect 1069 2124 1075 2136
rect 1053 1903 1059 1916
rect 1053 1897 1068 1903
rect 1085 1884 1091 2197
rect 1133 2124 1139 2136
rect 1197 2124 1203 2376
rect 1229 2324 1235 2456
rect 1245 2404 1251 2476
rect 1229 2304 1235 2316
rect 1213 2144 1219 2176
rect 1245 2124 1251 2356
rect 1261 2064 1267 2857
rect 1293 2784 1299 2796
rect 1309 2763 1315 2916
rect 1341 2904 1347 3077
rect 1501 3064 1507 3136
rect 1357 2964 1363 2996
rect 1501 2984 1507 3016
rect 1517 2984 1523 3036
rect 1533 2963 1539 3056
rect 1517 2957 1539 2963
rect 1373 2943 1379 2956
rect 1357 2937 1379 2943
rect 1293 2757 1315 2763
rect 1325 2897 1340 2903
rect 1293 2564 1299 2757
rect 1325 2664 1331 2897
rect 1309 2644 1315 2656
rect 1309 2544 1315 2636
rect 1341 2584 1347 2756
rect 1277 2323 1283 2536
rect 1277 2317 1299 2323
rect 1293 2284 1299 2317
rect 1309 2304 1315 2496
rect 1293 2264 1299 2276
rect 1309 2244 1315 2256
rect 1133 2024 1139 2036
rect 1117 1884 1123 1916
rect 1213 1904 1219 1936
rect 1229 1924 1235 2036
rect 1277 1983 1283 2156
rect 1309 2124 1315 2236
rect 1293 2004 1299 2036
rect 1277 1977 1299 1983
rect 1277 1904 1283 1956
rect 1293 1883 1299 1977
rect 1309 1964 1315 2056
rect 1325 2044 1331 2556
rect 1341 2304 1347 2436
rect 1357 2243 1363 2937
rect 1469 2924 1475 2936
rect 1373 2784 1379 2876
rect 1389 2704 1395 2916
rect 1434 2814 1446 2816
rect 1419 2806 1421 2814
rect 1429 2806 1431 2814
rect 1439 2806 1441 2814
rect 1449 2806 1451 2814
rect 1459 2806 1461 2814
rect 1434 2804 1446 2806
rect 1517 2784 1523 2957
rect 1565 2944 1571 3156
rect 1581 3004 1587 3096
rect 1613 2924 1619 3176
rect 1821 3144 1827 3336
rect 1853 3324 1859 3636
rect 1869 3584 1875 3676
rect 1885 3584 1891 3716
rect 1901 3484 1907 3556
rect 2077 3543 2083 3676
rect 2061 3537 2083 3543
rect 2045 3504 2051 3516
rect 1917 3404 1923 3496
rect 2061 3484 2067 3537
rect 1997 3424 2003 3456
rect 2013 3424 2019 3456
rect 1885 3364 1891 3376
rect 2013 3324 2019 3336
rect 1917 3284 1923 3296
rect 1837 3184 1843 3196
rect 1853 3163 1859 3236
rect 1933 3204 1939 3316
rect 1965 3284 1971 3316
rect 2029 3304 2035 3436
rect 2077 3324 2083 3376
rect 2093 3324 2099 4236
rect 2157 4184 2163 4256
rect 2189 4144 2195 4156
rect 2109 3764 2115 3956
rect 2205 3884 2211 4276
rect 2221 4184 2227 4236
rect 2253 4204 2259 4296
rect 2301 4184 2307 4316
rect 2317 4264 2323 4296
rect 2365 4284 2371 4376
rect 2429 4304 2435 4436
rect 2477 4324 2483 4436
rect 2525 4343 2531 4636
rect 2557 4604 2563 4856
rect 2573 4844 2579 4936
rect 2605 4864 2611 4956
rect 2621 4944 2627 4976
rect 2685 4964 2691 5296
rect 2621 4864 2627 4936
rect 2717 4924 2723 5094
rect 2749 5084 2755 5336
rect 2781 5224 2787 5316
rect 2781 5124 2787 5196
rect 2781 4924 2787 5016
rect 2797 4924 2803 5156
rect 2829 5104 2835 5316
rect 2845 4924 2851 5096
rect 2605 4784 2611 4816
rect 2701 4804 2707 4916
rect 2781 4904 2787 4916
rect 2701 4764 2707 4796
rect 2596 4717 2611 4723
rect 2573 4704 2579 4716
rect 2605 4584 2611 4717
rect 2589 4544 2595 4576
rect 2621 4564 2627 4616
rect 2637 4543 2643 4696
rect 2685 4664 2691 4696
rect 2701 4663 2707 4716
rect 2733 4684 2739 4836
rect 2701 4657 2716 4663
rect 2653 4584 2659 4656
rect 2733 4624 2739 4636
rect 2685 4584 2691 4596
rect 2669 4544 2675 4576
rect 2749 4564 2755 4836
rect 2861 4784 2867 5096
rect 2877 4943 2883 5076
rect 2893 5024 2899 5096
rect 2938 5014 2950 5016
rect 2923 5006 2925 5014
rect 2933 5006 2935 5014
rect 2943 5006 2945 5014
rect 2953 5006 2955 5014
rect 2963 5006 2965 5014
rect 2938 5004 2950 5006
rect 2989 4984 2995 5216
rect 3005 5184 3011 5457
rect 3437 5424 3443 5463
rect 3469 5404 3475 5463
rect 3501 5424 3507 5463
rect 3565 5404 3571 5463
rect 3597 5457 3619 5463
rect 3069 5326 3075 5356
rect 3213 5324 3219 5336
rect 3133 5164 3139 5236
rect 3053 5124 3059 5136
rect 3213 5124 3219 5316
rect 3261 5243 3267 5318
rect 3325 5304 3331 5336
rect 3341 5324 3347 5336
rect 3357 5243 3363 5376
rect 3437 5323 3443 5396
rect 3453 5344 3459 5376
rect 3469 5324 3475 5336
rect 3421 5317 3443 5323
rect 3421 5244 3427 5317
rect 3453 5284 3459 5316
rect 3261 5237 3283 5243
rect 3037 5004 3043 5096
rect 3101 4944 3107 4996
rect 2877 4937 2892 4943
rect 2845 4704 2851 4736
rect 2765 4584 2771 4696
rect 2829 4684 2835 4696
rect 2781 4664 2787 4676
rect 2877 4604 2883 4696
rect 2740 4557 2748 4563
rect 2781 4544 2787 4576
rect 2621 4537 2643 4543
rect 2621 4464 2627 4537
rect 2765 4524 2771 4536
rect 2829 4524 2835 4536
rect 2637 4504 2643 4516
rect 2717 4504 2723 4516
rect 2509 4337 2531 4343
rect 2509 4324 2515 4337
rect 2253 4164 2259 4176
rect 2349 4124 2355 4136
rect 2237 4104 2243 4116
rect 2285 4104 2291 4116
rect 2381 4084 2387 4136
rect 2397 4124 2403 4296
rect 2413 4224 2419 4296
rect 2429 4244 2435 4276
rect 2461 4264 2467 4276
rect 2285 3904 2291 3936
rect 2365 3904 2371 3936
rect 2381 3903 2387 4036
rect 2445 3924 2451 4236
rect 2461 4184 2467 4236
rect 2477 4224 2483 4276
rect 2525 4244 2531 4316
rect 2461 4144 2467 4156
rect 2477 4144 2483 4176
rect 2477 4084 2483 4116
rect 2381 3897 2403 3903
rect 2397 3884 2403 3897
rect 2493 3884 2499 4236
rect 2525 4144 2531 4156
rect 2541 4124 2547 4316
rect 2557 4144 2563 4396
rect 2605 4384 2611 4436
rect 2628 4337 2643 4343
rect 2573 4204 2579 4276
rect 2589 4244 2595 4316
rect 2637 4184 2643 4337
rect 2685 4284 2691 4316
rect 2701 4304 2707 4396
rect 2717 4317 2732 4323
rect 2717 4184 2723 4317
rect 2733 4204 2739 4236
rect 2509 4004 2515 4116
rect 2509 3884 2515 3936
rect 2557 3904 2563 4136
rect 2605 4064 2611 4096
rect 2621 3904 2627 3916
rect 2125 3704 2131 3836
rect 2141 3724 2147 3736
rect 2157 3724 2163 3836
rect 2205 3804 2211 3876
rect 2317 3864 2323 3876
rect 2269 3804 2275 3836
rect 2173 3764 2179 3796
rect 2205 3744 2211 3756
rect 2205 3664 2211 3716
rect 2109 3504 2115 3656
rect 1997 3284 2003 3296
rect 1949 3184 1955 3256
rect 1853 3157 1875 3163
rect 1645 3044 1651 3096
rect 1661 2944 1667 2956
rect 1677 2924 1683 2936
rect 1693 2924 1699 3096
rect 1709 3044 1715 3096
rect 1725 3024 1731 3136
rect 1773 3044 1779 3096
rect 1709 2944 1715 2956
rect 1741 2924 1747 2936
rect 1757 2924 1763 2956
rect 1597 2824 1603 2896
rect 1405 2523 1411 2656
rect 1437 2584 1443 2676
rect 1396 2517 1411 2523
rect 1421 2464 1427 2556
rect 1437 2464 1443 2496
rect 1434 2414 1446 2416
rect 1419 2406 1421 2414
rect 1429 2406 1431 2414
rect 1439 2406 1441 2414
rect 1449 2406 1451 2414
rect 1459 2406 1461 2414
rect 1434 2404 1446 2406
rect 1341 2237 1363 2243
rect 1341 2164 1347 2237
rect 1469 2224 1475 2296
rect 1357 2144 1363 2176
rect 1405 2144 1411 2156
rect 1421 2124 1427 2156
rect 1341 1964 1347 2036
rect 1434 2014 1446 2016
rect 1419 2006 1421 2014
rect 1429 2006 1431 2014
rect 1439 2006 1441 2014
rect 1449 2006 1451 2014
rect 1459 2006 1461 2014
rect 1434 2004 1446 2006
rect 1373 1984 1379 1996
rect 1309 1904 1315 1936
rect 1341 1904 1347 1916
rect 1325 1884 1331 1896
rect 1069 1784 1075 1856
rect 781 1724 787 1736
rect 756 1717 771 1723
rect 765 1584 771 1717
rect 781 1544 787 1576
rect 749 1524 755 1536
rect 813 1503 819 1716
rect 797 1497 819 1503
rect 829 1517 844 1523
rect 749 1384 755 1456
rect 797 1424 803 1497
rect 829 1464 835 1517
rect 861 1484 867 1736
rect 877 1524 883 1756
rect 733 1364 739 1376
rect 637 1344 643 1356
rect 701 1344 707 1356
rect 797 1344 803 1416
rect 861 1404 867 1436
rect 877 1384 883 1476
rect 893 1463 899 1496
rect 909 1484 915 1736
rect 925 1544 931 1716
rect 925 1504 931 1516
rect 893 1457 924 1463
rect 941 1384 947 1656
rect 669 1284 675 1296
rect 269 1064 275 1096
rect 285 1084 291 1276
rect 605 1264 611 1276
rect 301 1043 307 1256
rect 477 1104 483 1236
rect 493 1104 499 1116
rect 749 1104 755 1336
rect 893 1324 899 1336
rect 909 1324 915 1336
rect 797 1224 803 1316
rect 893 1304 899 1316
rect 829 1104 835 1276
rect 845 1124 851 1136
rect 909 1104 915 1316
rect 941 1124 947 1316
rect 957 1144 963 1456
rect 1005 1384 1011 1716
rect 1037 1504 1043 1736
rect 1085 1724 1091 1756
rect 1085 1584 1091 1696
rect 1069 1544 1075 1576
rect 1101 1524 1107 1536
rect 1069 1483 1075 1516
rect 1069 1477 1091 1483
rect 1037 1464 1043 1476
rect 1069 1364 1075 1456
rect 1085 1384 1091 1477
rect 1101 1344 1107 1436
rect 1117 1343 1123 1776
rect 1133 1704 1139 1880
rect 1277 1877 1299 1883
rect 1181 1724 1187 1736
rect 1229 1544 1235 1836
rect 1245 1764 1251 1796
rect 1261 1743 1267 1756
rect 1252 1737 1267 1743
rect 1165 1444 1171 1464
rect 1213 1444 1219 1476
rect 1229 1464 1235 1476
rect 1181 1364 1187 1436
rect 1261 1364 1267 1436
rect 1117 1337 1132 1343
rect 1021 1184 1027 1196
rect 1053 1164 1059 1336
rect 1133 1324 1139 1336
rect 1117 1303 1123 1316
rect 1149 1303 1155 1356
rect 1261 1324 1267 1356
rect 1117 1297 1155 1303
rect 1181 1264 1187 1316
rect 957 1104 963 1116
rect 301 1037 316 1043
rect 237 1017 259 1023
rect 237 984 243 1017
rect 157 944 163 976
rect 285 944 291 1036
rect 13 884 19 896
rect 45 884 51 916
rect 13 784 19 856
rect 13 564 19 656
rect 45 564 51 876
rect 61 864 67 936
rect 61 684 67 696
rect 141 684 147 736
rect 157 724 163 936
rect 173 724 179 936
rect 237 784 243 916
rect 157 704 163 716
rect 77 664 83 676
rect 173 663 179 716
rect 189 684 195 696
rect 164 657 179 663
rect 77 564 83 636
rect 109 584 115 636
rect 157 584 163 656
rect 29 523 35 556
rect 45 544 51 556
rect 20 517 35 523
rect 205 504 211 676
rect 237 624 243 656
rect 253 644 259 656
rect 237 524 243 576
rect 269 543 275 936
rect 317 924 323 1036
rect 365 1024 371 1096
rect 381 943 387 1056
rect 397 964 403 1056
rect 372 937 387 943
rect 445 924 451 1096
rect 365 884 371 896
rect 285 723 291 736
rect 349 724 355 836
rect 285 717 307 723
rect 301 704 307 717
rect 365 704 371 876
rect 461 864 467 1036
rect 477 964 483 1076
rect 509 1064 515 1076
rect 557 1064 563 1096
rect 461 743 467 836
rect 445 737 467 743
rect 445 703 451 737
rect 445 697 467 703
rect 285 684 291 696
rect 461 684 467 697
rect 477 684 483 696
rect 493 684 499 856
rect 436 677 451 683
rect 301 664 307 676
rect 285 544 291 556
rect 365 544 371 556
rect 260 537 275 543
rect 253 503 259 536
rect 301 504 307 516
rect 333 504 339 516
rect 253 497 275 503
rect 45 384 51 496
rect 141 384 147 496
rect 109 284 115 296
rect 125 263 131 276
rect 109 257 131 263
rect 109 244 115 257
rect 61 184 67 236
rect 125 184 131 236
rect 141 184 147 296
rect 189 284 195 316
rect 221 284 227 316
rect 269 304 275 497
rect 349 304 355 536
rect 397 344 403 636
rect 445 564 451 677
rect 477 644 483 676
rect 509 563 515 1036
rect 525 984 531 1036
rect 541 964 547 1056
rect 557 904 563 1016
rect 573 964 579 1056
rect 589 964 595 1056
rect 653 964 659 1056
rect 701 984 707 1076
rect 733 964 739 1056
rect 621 944 627 956
rect 637 903 643 916
rect 685 903 691 956
rect 637 897 691 903
rect 541 724 547 736
rect 557 583 563 896
rect 749 703 755 1096
rect 829 1044 835 1096
rect 797 1024 803 1036
rect 765 964 771 1016
rect 877 1004 883 1096
rect 909 1084 915 1096
rect 893 1063 899 1076
rect 973 1063 979 1136
rect 989 1064 995 1096
rect 1021 1084 1027 1116
rect 1149 1104 1155 1116
rect 893 1057 915 1063
rect 797 984 803 996
rect 909 984 915 1057
rect 957 1057 979 1063
rect 781 904 787 956
rect 813 944 819 976
rect 861 924 867 956
rect 877 904 883 976
rect 925 963 931 1036
rect 957 964 963 1057
rect 1053 1024 1059 1076
rect 1069 1003 1075 1096
rect 1165 1044 1171 1096
rect 1101 1024 1107 1036
rect 1053 997 1075 1003
rect 909 957 931 963
rect 845 844 851 876
rect 861 864 867 876
rect 749 697 764 703
rect 573 677 588 683
rect 573 584 579 677
rect 493 557 515 563
rect 541 577 563 583
rect 493 524 499 557
rect 509 444 515 536
rect 541 524 547 577
rect 669 564 675 656
rect 685 644 691 696
rect 813 683 819 716
rect 852 697 876 703
rect 909 684 915 957
rect 941 944 947 956
rect 1037 944 1043 956
rect 1053 944 1059 997
rect 925 924 931 936
rect 957 924 963 936
rect 1012 897 1027 903
rect 804 677 819 683
rect 701 604 707 676
rect 749 564 755 656
rect 781 564 787 636
rect 749 544 755 556
rect 797 544 803 656
rect 813 644 819 677
rect 845 664 851 676
rect 845 584 851 596
rect 861 544 867 556
rect 909 544 915 556
rect 589 524 595 536
rect 925 523 931 796
rect 941 784 947 836
rect 1021 784 1027 897
rect 957 704 963 716
rect 1005 684 1011 696
rect 909 517 931 523
rect 653 504 659 516
rect 669 504 675 516
rect 845 504 851 516
rect 397 304 403 336
rect 429 304 435 316
rect 189 244 195 276
rect 189 184 195 196
rect 13 144 19 156
rect 45 144 51 156
rect 205 104 211 236
rect 221 204 227 276
rect 253 140 259 256
rect 285 184 291 296
rect 301 244 307 296
rect 349 264 355 296
rect 461 284 467 436
rect 509 284 515 436
rect 468 277 476 283
rect 397 264 403 276
rect 317 144 323 256
rect 333 204 339 256
rect 333 164 339 196
rect 285 104 291 136
rect 381 124 387 236
rect 461 184 467 216
rect 509 184 515 276
rect 413 164 419 176
rect 509 144 515 156
rect 525 124 531 256
rect 541 124 547 296
rect 605 284 611 296
rect 653 244 659 276
rect 669 264 675 336
rect 685 304 691 316
rect 701 263 707 276
rect 701 257 716 263
rect 605 164 611 196
rect 621 184 627 236
rect 637 184 643 216
rect 669 184 675 236
rect 733 164 739 236
rect 749 164 755 356
rect 781 264 787 376
rect 813 224 819 316
rect 845 304 851 316
rect 909 303 915 517
rect 925 364 931 436
rect 941 384 947 556
rect 957 524 963 676
rect 1021 584 1027 756
rect 1053 684 1059 936
rect 1085 664 1091 676
rect 989 564 995 576
rect 1005 544 1011 556
rect 1037 524 1043 536
rect 1053 484 1059 516
rect 1069 384 1075 656
rect 1085 584 1091 656
rect 1101 584 1107 996
rect 1181 924 1187 1256
rect 1213 1244 1219 1296
rect 1277 1244 1283 1877
rect 1357 1864 1363 1976
rect 1373 1944 1379 1976
rect 1389 1904 1395 1956
rect 1485 1924 1491 2636
rect 1501 2584 1507 2696
rect 1517 2504 1523 2536
rect 1533 2444 1539 2796
rect 1549 2584 1555 2696
rect 1613 2684 1619 2876
rect 1645 2764 1651 2916
rect 1693 2904 1699 2916
rect 1789 2884 1795 3136
rect 1805 2924 1811 3036
rect 1821 3004 1827 3116
rect 1837 3044 1843 3096
rect 1853 2984 1859 3116
rect 1869 3044 1875 3157
rect 1949 3144 1955 3156
rect 1949 3104 1955 3136
rect 1885 3084 1891 3096
rect 1869 2944 1875 2976
rect 1821 2904 1827 2916
rect 1549 2544 1555 2556
rect 1565 2384 1571 2536
rect 1581 2464 1587 2556
rect 1597 2544 1603 2680
rect 1661 2664 1667 2756
rect 1677 2704 1683 2776
rect 1741 2744 1747 2836
rect 1709 2724 1715 2736
rect 1773 2724 1779 2776
rect 1869 2764 1875 2896
rect 1684 2677 1699 2683
rect 1636 2657 1651 2663
rect 1629 2504 1635 2556
rect 1645 2483 1651 2657
rect 1629 2477 1651 2483
rect 1517 2124 1523 2356
rect 1613 2344 1619 2436
rect 1629 2384 1635 2477
rect 1533 2244 1539 2336
rect 1661 2324 1667 2656
rect 1693 2584 1699 2677
rect 1789 2624 1795 2696
rect 1837 2664 1843 2696
rect 1837 2584 1843 2656
rect 1853 2644 1859 2656
rect 1725 2524 1731 2556
rect 1757 2544 1763 2556
rect 1741 2523 1747 2536
rect 1885 2524 1891 3076
rect 1965 3064 1971 3136
rect 1933 2884 1939 3056
rect 1981 3024 1987 3236
rect 2013 3184 2019 3216
rect 1997 3064 2003 3096
rect 1917 2784 1923 2836
rect 1949 2824 1955 2916
rect 1965 2904 1971 2956
rect 2013 2944 2019 3076
rect 2029 2984 2035 3276
rect 2045 2944 2051 2956
rect 2045 2924 2051 2936
rect 2061 2924 2067 3096
rect 1981 2883 1987 2916
rect 1965 2877 1987 2883
rect 1741 2517 1763 2523
rect 1613 2297 1628 2303
rect 1517 2084 1523 2096
rect 1533 2063 1539 2116
rect 1565 2084 1571 2296
rect 1517 2057 1539 2063
rect 1517 1944 1523 2057
rect 1565 1984 1571 2056
rect 1549 1944 1555 1976
rect 1581 1964 1587 2116
rect 1597 2084 1603 2096
rect 1613 2064 1619 2297
rect 1645 2303 1651 2316
rect 1645 2297 1660 2303
rect 1629 2144 1635 2176
rect 1597 1984 1603 2016
rect 1293 1784 1299 1796
rect 1357 1764 1363 1796
rect 1373 1784 1379 1896
rect 1293 1704 1299 1716
rect 1309 1703 1315 1756
rect 1325 1724 1331 1756
rect 1341 1744 1347 1756
rect 1389 1724 1395 1796
rect 1405 1764 1411 1916
rect 1565 1904 1571 1956
rect 1613 1944 1619 1956
rect 1517 1804 1523 1876
rect 1501 1783 1507 1796
rect 1501 1777 1516 1783
rect 1581 1764 1587 1916
rect 1629 1904 1635 2076
rect 1645 2024 1651 2116
rect 1629 1764 1635 1776
rect 1549 1724 1555 1736
rect 1309 1697 1436 1703
rect 1533 1703 1539 1716
rect 1492 1697 1539 1703
rect 1357 1584 1363 1676
rect 1434 1614 1446 1616
rect 1419 1606 1421 1614
rect 1429 1606 1431 1614
rect 1439 1606 1441 1614
rect 1449 1606 1451 1614
rect 1459 1606 1461 1614
rect 1434 1604 1446 1606
rect 1485 1584 1491 1636
rect 1293 1324 1299 1376
rect 1309 1324 1315 1496
rect 1357 1457 1372 1463
rect 1341 1444 1347 1456
rect 1341 1364 1347 1396
rect 1197 944 1203 1036
rect 1213 924 1219 1216
rect 1229 1064 1235 1076
rect 1245 1064 1251 1236
rect 1357 1204 1363 1457
rect 1373 1324 1379 1336
rect 1389 1244 1395 1496
rect 1501 1484 1507 1676
rect 1565 1584 1571 1736
rect 1661 1724 1667 2276
rect 1677 2104 1683 2436
rect 1725 2284 1731 2516
rect 1741 2384 1747 2436
rect 1757 2384 1763 2517
rect 1693 2244 1699 2276
rect 1741 2264 1747 2296
rect 1757 2264 1763 2376
rect 1677 2084 1683 2096
rect 1693 2063 1699 2096
rect 1684 2057 1699 2063
rect 1677 1944 1683 1956
rect 1709 1943 1715 2036
rect 1725 1964 1731 2116
rect 1709 1937 1731 1943
rect 1677 1724 1683 1736
rect 1581 1664 1587 1716
rect 1661 1644 1667 1716
rect 1693 1684 1699 1716
rect 1709 1664 1715 1916
rect 1725 1884 1731 1937
rect 1741 1884 1747 1896
rect 1757 1664 1763 2256
rect 1789 2184 1795 2336
rect 1853 2264 1859 2516
rect 1885 2404 1891 2476
rect 1901 2384 1907 2516
rect 1917 2503 1923 2636
rect 1949 2563 1955 2756
rect 1965 2724 1971 2877
rect 2013 2704 2019 2836
rect 2045 2704 2051 2856
rect 1965 2624 1971 2656
rect 1949 2557 1971 2563
rect 1965 2524 1971 2557
rect 1981 2544 1987 2556
rect 1997 2524 2003 2656
rect 2029 2564 2035 2676
rect 2045 2524 2051 2616
rect 1917 2497 1939 2503
rect 1933 2364 1939 2497
rect 1869 2284 1875 2296
rect 1901 2184 1907 2276
rect 1933 2203 1939 2356
rect 1965 2344 1971 2516
rect 1997 2324 2003 2516
rect 2029 2484 2035 2496
rect 2061 2484 2067 2636
rect 2077 2543 2083 3216
rect 2093 3184 2099 3296
rect 2109 3224 2115 3496
rect 2141 3304 2147 3636
rect 2180 3517 2195 3523
rect 2157 3424 2163 3456
rect 2189 3444 2195 3517
rect 2221 3484 2227 3796
rect 2269 3764 2275 3776
rect 2253 3744 2259 3756
rect 2317 3744 2323 3796
rect 2333 3744 2339 3836
rect 2413 3764 2419 3796
rect 2237 3504 2243 3716
rect 2301 3564 2307 3636
rect 2253 3504 2259 3536
rect 2301 3444 2307 3516
rect 2333 3504 2339 3716
rect 2365 3664 2371 3716
rect 2397 3504 2403 3656
rect 2349 3464 2355 3476
rect 2141 3184 2147 3196
rect 2157 3164 2163 3316
rect 2093 3104 2099 3116
rect 2093 2824 2099 3096
rect 2109 3064 2115 3136
rect 2125 3043 2131 3136
rect 2173 3104 2179 3436
rect 2237 3424 2243 3436
rect 2237 3364 2243 3396
rect 2285 3344 2291 3436
rect 2317 3343 2323 3436
rect 2429 3344 2435 3836
rect 2461 3744 2467 3816
rect 2493 3524 2499 3716
rect 2525 3684 2531 3716
rect 2573 3704 2579 3836
rect 2621 3744 2627 3836
rect 2637 3784 2643 4136
rect 2653 4124 2659 4136
rect 2669 4024 2675 4116
rect 2701 3923 2707 4176
rect 2749 4163 2755 4256
rect 2765 4184 2771 4516
rect 2797 4304 2803 4376
rect 2781 4224 2787 4236
rect 2749 4157 2771 4163
rect 2765 4144 2771 4157
rect 2797 4144 2803 4176
rect 2861 4164 2867 4556
rect 2893 4543 2899 4876
rect 2925 4864 2931 4896
rect 2989 4684 2995 4836
rect 3037 4804 3043 4916
rect 3053 4884 3059 4936
rect 2938 4614 2950 4616
rect 2923 4606 2925 4614
rect 2933 4606 2935 4614
rect 2943 4606 2945 4614
rect 2953 4606 2955 4614
rect 2963 4606 2965 4614
rect 2938 4604 2950 4606
rect 2893 4537 2915 4543
rect 2909 4444 2915 4537
rect 2925 4524 2931 4536
rect 2909 4283 2915 4336
rect 2989 4304 2995 4616
rect 3021 4544 3027 4556
rect 3012 4517 3027 4523
rect 3005 4304 3011 4496
rect 3021 4384 3027 4517
rect 3053 4504 3059 4876
rect 3085 4844 3091 4916
rect 3069 4684 3075 4696
rect 3085 4624 3091 4636
rect 3117 4544 3123 5096
rect 3133 4884 3139 4936
rect 3149 4704 3155 5096
rect 3213 5084 3219 5116
rect 3245 5104 3251 5136
rect 3181 4944 3187 5056
rect 3229 4904 3235 5016
rect 3261 4903 3267 5136
rect 3277 5004 3283 5237
rect 3341 5237 3363 5243
rect 3309 5104 3315 5116
rect 3293 4944 3299 4956
rect 3277 4924 3283 4936
rect 3261 4897 3283 4903
rect 3165 4884 3171 4896
rect 3165 4784 3171 4836
rect 3261 4704 3267 4876
rect 3037 4484 3043 4496
rect 3053 4384 3059 4476
rect 2893 4277 2915 4283
rect 2893 4184 2899 4277
rect 2938 4214 2950 4216
rect 2923 4206 2925 4214
rect 2933 4206 2935 4214
rect 2943 4206 2945 4214
rect 2953 4206 2955 4214
rect 2963 4206 2965 4214
rect 2938 4204 2950 4206
rect 2733 4024 2739 4136
rect 2781 4124 2787 4136
rect 2845 4084 2851 4156
rect 2909 4144 2915 4176
rect 2701 3917 2716 3923
rect 2701 3904 2707 3917
rect 2733 3863 2739 3996
rect 2765 3884 2771 4076
rect 2845 4004 2851 4076
rect 2877 3924 2883 4016
rect 2717 3857 2739 3863
rect 2669 3804 2675 3836
rect 2717 3744 2723 3857
rect 2605 3724 2611 3736
rect 2733 3724 2739 3836
rect 2781 3824 2787 3836
rect 2781 3744 2787 3796
rect 2797 3724 2803 3916
rect 2845 3884 2851 3896
rect 2877 3884 2883 3916
rect 2925 3884 2931 4156
rect 2989 4124 2995 4236
rect 3021 4184 3027 4376
rect 3037 4124 3043 4236
rect 3021 4117 3036 4123
rect 2989 4104 2995 4116
rect 2989 3964 2995 4096
rect 2861 3864 2867 3876
rect 2861 3764 2867 3856
rect 2877 3804 2883 3836
rect 2938 3814 2950 3816
rect 2923 3806 2925 3814
rect 2933 3806 2935 3814
rect 2943 3806 2945 3814
rect 2953 3806 2955 3814
rect 2963 3806 2965 3814
rect 2938 3804 2950 3806
rect 3005 3764 3011 3836
rect 2445 3424 2451 3456
rect 2461 3384 2467 3436
rect 2317 3337 2339 3343
rect 2196 3317 2211 3323
rect 2205 3284 2211 3317
rect 2109 3037 2131 3043
rect 2109 2984 2115 3037
rect 2109 2704 2115 2936
rect 2125 2924 2131 2956
rect 2141 2944 2147 2976
rect 2141 2903 2147 2916
rect 2189 2904 2195 2976
rect 2125 2897 2147 2903
rect 2093 2624 2099 2656
rect 2109 2644 2115 2676
rect 2125 2604 2131 2897
rect 2205 2864 2211 3276
rect 2317 3224 2323 3316
rect 2301 3144 2307 3156
rect 2221 3064 2227 3136
rect 2237 3104 2243 3116
rect 2285 3064 2291 3136
rect 2333 3124 2339 3337
rect 2349 3324 2355 3336
rect 2301 3104 2307 3116
rect 2269 2964 2275 2996
rect 2237 2944 2243 2956
rect 2301 2944 2307 2956
rect 2301 2864 2307 2916
rect 2077 2537 2099 2543
rect 1972 2317 1987 2323
rect 1933 2197 1955 2203
rect 1773 2084 1779 2156
rect 1789 2124 1795 2176
rect 1853 2124 1859 2176
rect 1949 2124 1955 2197
rect 1853 2083 1859 2096
rect 1853 2077 1900 2083
rect 1805 1984 1811 2076
rect 1837 1984 1843 2076
rect 1917 2064 1923 2116
rect 1965 2104 1971 2236
rect 1917 1984 1923 2016
rect 1837 1944 1843 1976
rect 1853 1904 1859 1956
rect 1901 1944 1907 1976
rect 1869 1884 1875 1916
rect 1917 1904 1923 1956
rect 1981 1924 1987 2317
rect 1997 2244 2003 2276
rect 2013 2143 2019 2456
rect 2029 2164 2035 2336
rect 2045 2324 2051 2356
rect 2045 2284 2051 2296
rect 2077 2283 2083 2436
rect 2093 2304 2099 2537
rect 2141 2504 2147 2636
rect 2157 2624 2163 2656
rect 2189 2644 2195 2676
rect 2157 2523 2163 2596
rect 2173 2543 2179 2636
rect 2205 2624 2211 2836
rect 2285 2704 2291 2856
rect 2173 2537 2188 2543
rect 2157 2517 2172 2523
rect 2221 2504 2227 2636
rect 2237 2624 2243 2656
rect 2237 2524 2243 2536
rect 2253 2524 2259 2556
rect 2269 2544 2275 2696
rect 2285 2564 2291 2636
rect 2317 2603 2323 3096
rect 2333 2844 2339 2916
rect 2365 2904 2371 3296
rect 2397 3004 2403 3336
rect 2445 3244 2451 3276
rect 2445 3144 2451 3156
rect 2413 3124 2419 3136
rect 2477 3124 2483 3416
rect 2509 3304 2515 3316
rect 2525 3304 2531 3556
rect 2589 3504 2595 3636
rect 2557 3343 2563 3496
rect 2621 3484 2627 3716
rect 2605 3477 2620 3483
rect 2605 3463 2611 3477
rect 2596 3457 2611 3463
rect 2557 3337 2579 3343
rect 2493 3264 2499 3276
rect 2429 3104 2435 3116
rect 2381 2964 2387 2996
rect 2333 2704 2339 2836
rect 2397 2724 2403 2896
rect 2413 2824 2419 3096
rect 2429 2944 2435 2996
rect 2477 2984 2483 3096
rect 2509 3083 2515 3236
rect 2541 3164 2547 3316
rect 2541 3084 2547 3096
rect 2509 3077 2531 3083
rect 2509 3044 2515 3056
rect 2525 3044 2531 3077
rect 2445 2944 2451 2976
rect 2493 2964 2499 2996
rect 2541 2984 2547 3056
rect 2557 2984 2563 3036
rect 2333 2624 2339 2696
rect 2365 2624 2371 2656
rect 2413 2644 2419 2676
rect 2461 2644 2467 2716
rect 2477 2684 2483 2876
rect 2317 2597 2339 2603
rect 2317 2544 2323 2576
rect 2237 2484 2243 2516
rect 2269 2464 2275 2536
rect 2333 2523 2339 2597
rect 2365 2524 2371 2596
rect 2381 2544 2387 2636
rect 2324 2517 2339 2523
rect 2125 2343 2131 2436
rect 2125 2337 2147 2343
rect 2141 2323 2147 2337
rect 2141 2317 2163 2323
rect 2125 2297 2140 2303
rect 2109 2284 2115 2296
rect 2077 2277 2099 2283
rect 2077 2184 2083 2256
rect 2093 2164 2099 2277
rect 2109 2184 2115 2256
rect 2004 2137 2019 2143
rect 2045 2124 2051 2136
rect 2029 2044 2035 2096
rect 2061 2064 2067 2076
rect 2109 2004 2115 2036
rect 2125 1944 2131 2297
rect 2141 2084 2147 2176
rect 2157 2124 2163 2317
rect 2189 2264 2195 2296
rect 2205 2284 2211 2456
rect 2269 2344 2275 2436
rect 2301 2284 2307 2336
rect 2317 2304 2323 2516
rect 2349 2304 2355 2516
rect 2397 2304 2403 2616
rect 2413 2564 2419 2596
rect 2445 2504 2451 2636
rect 2493 2584 2499 2676
rect 2509 2604 2515 2876
rect 2541 2864 2547 2916
rect 2557 2704 2563 2716
rect 2573 2684 2579 3337
rect 2605 3343 2611 3436
rect 2621 3424 2627 3456
rect 2621 3344 2627 3356
rect 2637 3344 2643 3636
rect 2685 3504 2691 3636
rect 2733 3504 2739 3536
rect 2701 3344 2707 3436
rect 2596 3337 2611 3343
rect 2605 3184 2611 3316
rect 2637 3284 2643 3316
rect 2605 3043 2611 3176
rect 2637 3144 2643 3276
rect 2637 3104 2643 3116
rect 2669 3104 2675 3216
rect 2589 3037 2611 3043
rect 2589 2924 2595 3037
rect 2621 2964 2627 2996
rect 2669 2984 2675 3076
rect 2637 2944 2643 2976
rect 2589 2844 2595 2916
rect 2653 2724 2659 2756
rect 2669 2744 2675 2756
rect 2509 2524 2515 2596
rect 2253 2244 2259 2276
rect 2429 2264 2435 2276
rect 2173 2064 2179 2096
rect 2221 2084 2227 2236
rect 2269 2124 2275 2236
rect 2317 2224 2323 2256
rect 1789 1824 1795 1856
rect 1853 1824 1859 1836
rect 1837 1784 1843 1796
rect 1789 1724 1795 1756
rect 1885 1724 1891 1736
rect 1821 1684 1827 1716
rect 1869 1703 1875 1716
rect 1869 1697 1891 1703
rect 1869 1684 1875 1697
rect 1885 1684 1891 1697
rect 1677 1584 1683 1656
rect 1597 1504 1603 1516
rect 1405 1304 1411 1356
rect 1389 1224 1395 1236
rect 1485 1224 1491 1456
rect 1517 1444 1523 1496
rect 1533 1423 1539 1456
rect 1549 1444 1555 1476
rect 1517 1417 1539 1423
rect 1517 1384 1523 1417
rect 1549 1364 1555 1436
rect 1565 1384 1571 1476
rect 1613 1464 1619 1476
rect 1581 1417 1619 1423
rect 1581 1404 1587 1417
rect 1597 1364 1603 1396
rect 1613 1364 1619 1417
rect 1709 1384 1715 1636
rect 1901 1624 1907 1876
rect 1917 1584 1923 1676
rect 1933 1644 1939 1916
rect 1997 1903 2003 1916
rect 2077 1904 2083 1936
rect 1997 1897 2012 1903
rect 2109 1903 2115 1916
rect 2157 1904 2163 2036
rect 2189 1984 2195 2016
rect 2205 1904 2211 2036
rect 2237 1984 2243 2056
rect 2269 1917 2284 1923
rect 2269 1904 2275 1917
rect 2109 1897 2124 1903
rect 1981 1884 1987 1896
rect 1949 1744 1955 1836
rect 1965 1804 1971 1856
rect 2045 1844 2051 1876
rect 2045 1764 2051 1796
rect 1949 1623 1955 1716
rect 2045 1684 2051 1736
rect 2061 1724 2067 1836
rect 2093 1824 2099 1896
rect 2157 1844 2163 1876
rect 2109 1784 2115 1816
rect 2157 1764 2163 1796
rect 2221 1784 2227 1856
rect 2237 1824 2243 1896
rect 2253 1744 2259 1896
rect 2269 1764 2275 1796
rect 2061 1704 2067 1716
rect 1949 1617 1971 1623
rect 1789 1504 1795 1516
rect 1789 1464 1795 1496
rect 1933 1484 1939 1496
rect 1828 1457 1843 1463
rect 1508 1337 1532 1343
rect 1549 1324 1555 1356
rect 1434 1214 1446 1216
rect 1419 1206 1421 1214
rect 1429 1206 1431 1214
rect 1439 1206 1441 1214
rect 1449 1206 1451 1214
rect 1459 1206 1461 1214
rect 1434 1204 1446 1206
rect 1309 1124 1315 1196
rect 1277 1064 1283 1076
rect 1309 964 1315 1036
rect 1341 1024 1347 1096
rect 1357 1063 1363 1076
rect 1357 1057 1372 1063
rect 1389 984 1395 1196
rect 1581 1184 1587 1356
rect 1597 1344 1603 1356
rect 1661 1344 1667 1376
rect 1837 1364 1843 1457
rect 1869 1364 1875 1476
rect 1933 1464 1939 1476
rect 1805 1324 1811 1336
rect 1613 1304 1619 1316
rect 1613 1224 1619 1236
rect 1405 1064 1411 1076
rect 1421 1044 1427 1096
rect 1533 1064 1539 1156
rect 1597 1103 1603 1196
rect 1588 1097 1603 1103
rect 1629 1084 1635 1296
rect 1645 1224 1651 1296
rect 1757 1184 1763 1316
rect 1780 1297 1795 1303
rect 1661 1104 1667 1136
rect 1773 1064 1779 1076
rect 1789 1064 1795 1297
rect 1837 1084 1843 1316
rect 1869 1304 1875 1356
rect 1901 1224 1907 1456
rect 1933 1383 1939 1456
rect 1917 1377 1939 1383
rect 1853 1084 1859 1116
rect 1172 917 1180 923
rect 1277 904 1283 936
rect 1309 924 1315 956
rect 1517 944 1523 1036
rect 1533 1024 1539 1056
rect 1613 1044 1619 1056
rect 1661 950 1667 1036
rect 1821 1024 1827 1076
rect 1677 984 1683 1016
rect 1837 1004 1843 1056
rect 1885 956 1891 1116
rect 1917 1084 1923 1377
rect 1933 1344 1939 1356
rect 1933 1184 1939 1336
rect 1949 1184 1955 1196
rect 1901 1004 1907 1056
rect 1933 1024 1939 1096
rect 1949 943 1955 1056
rect 1940 937 1955 943
rect 1133 764 1139 836
rect 1181 724 1187 836
rect 1229 723 1235 836
rect 1277 784 1283 836
rect 1325 804 1331 936
rect 1341 764 1347 936
rect 1437 924 1443 936
rect 1549 884 1555 916
rect 1389 784 1395 876
rect 1434 814 1446 816
rect 1419 806 1421 814
rect 1429 806 1431 814
rect 1439 806 1441 814
rect 1449 806 1451 814
rect 1459 806 1461 814
rect 1434 804 1446 806
rect 1213 717 1235 723
rect 1213 684 1219 717
rect 1229 684 1235 696
rect 1148 664 1156 670
rect 1181 564 1187 664
rect 1293 624 1299 636
rect 893 297 915 303
rect 893 184 899 297
rect 909 264 915 276
rect 909 184 915 256
rect 925 224 931 316
rect 877 164 883 176
rect 573 144 579 156
rect 605 144 611 156
rect 733 124 739 156
rect 749 144 755 156
rect 941 144 947 376
rect 957 304 963 316
rect 989 304 995 356
rect 1117 284 1123 336
rect 973 244 979 276
rect 1133 264 1139 296
rect 1021 244 1027 256
rect 1085 204 1091 256
rect 1165 244 1171 536
rect 1197 284 1203 436
rect 1213 304 1219 556
rect 1261 544 1267 556
rect 1309 504 1315 536
rect 1325 524 1331 716
rect 1341 704 1347 736
rect 1501 704 1507 716
rect 1517 704 1523 756
rect 1357 684 1363 696
rect 1341 664 1347 676
rect 1357 624 1363 676
rect 1357 584 1363 596
rect 1389 584 1395 656
rect 1485 564 1491 636
rect 1517 604 1523 696
rect 1549 684 1555 876
rect 1629 744 1635 936
rect 1613 704 1619 716
rect 1597 684 1603 696
rect 1629 684 1635 716
rect 1661 664 1667 736
rect 1565 584 1571 656
rect 1661 604 1667 656
rect 1533 544 1539 556
rect 1629 544 1635 596
rect 1645 544 1651 556
rect 1677 544 1683 636
rect 1277 324 1283 476
rect 1325 384 1331 516
rect 1341 484 1347 536
rect 1357 384 1363 496
rect 1389 364 1395 516
rect 1421 504 1427 536
rect 1469 464 1475 496
rect 1501 484 1507 516
rect 1434 414 1446 416
rect 1419 406 1421 414
rect 1429 406 1431 414
rect 1439 406 1441 414
rect 1449 406 1451 414
rect 1459 406 1461 414
rect 1434 404 1446 406
rect 1341 304 1347 356
rect 1405 304 1411 316
rect 1165 184 1171 236
rect 1005 164 1011 176
rect 1229 164 1235 256
rect 1021 144 1027 156
rect 1229 144 1235 156
rect 1245 144 1251 276
rect 1261 184 1267 296
rect 1293 244 1299 256
rect 1325 204 1331 296
rect 1341 184 1347 296
rect 1421 264 1427 276
rect 1309 164 1315 176
rect 1437 144 1443 216
rect 1517 184 1523 536
rect 1693 524 1699 696
rect 1725 664 1731 936
rect 1789 784 1795 896
rect 1821 884 1827 936
rect 1901 784 1907 876
rect 1949 744 1955 836
rect 1965 784 1971 1617
rect 1997 1363 2003 1636
rect 2013 1584 2019 1616
rect 2125 1584 2131 1656
rect 2157 1524 2163 1736
rect 2189 1704 2195 1716
rect 2061 1497 2076 1503
rect 2013 1384 2019 1396
rect 1997 1357 2019 1363
rect 1997 1324 2003 1336
rect 1981 1204 1987 1316
rect 2013 1184 2019 1357
rect 2029 1304 2035 1336
rect 2045 1304 2051 1356
rect 2061 1264 2067 1497
rect 2077 1324 2083 1356
rect 2093 1303 2099 1476
rect 2141 1344 2147 1456
rect 2157 1404 2163 1476
rect 2157 1364 2163 1396
rect 2173 1323 2179 1676
rect 2221 1584 2227 1696
rect 2253 1484 2259 1496
rect 2253 1383 2259 1476
rect 2237 1377 2259 1383
rect 2189 1344 2195 1356
rect 2189 1324 2195 1336
rect 2157 1317 2179 1323
rect 2077 1297 2099 1303
rect 2061 1224 2067 1256
rect 2077 1184 2083 1297
rect 2141 1184 2147 1316
rect 2052 1097 2067 1103
rect 1981 944 1987 1096
rect 2029 1083 2035 1096
rect 2029 1077 2051 1083
rect 2004 1057 2019 1063
rect 1997 964 2003 1016
rect 2013 984 2019 1057
rect 1981 924 1987 936
rect 1997 824 2003 956
rect 2029 924 2035 996
rect 2045 984 2051 1077
rect 2061 864 2067 1097
rect 2093 1044 2099 1076
rect 2125 1064 2131 1096
rect 2077 940 2083 996
rect 2093 963 2099 1036
rect 2157 984 2163 1317
rect 2189 1297 2204 1303
rect 2189 1204 2195 1297
rect 2221 1283 2227 1316
rect 2205 1277 2227 1283
rect 2205 1184 2211 1277
rect 2237 1243 2243 1377
rect 2253 1304 2259 1356
rect 2237 1237 2259 1243
rect 2253 1184 2259 1237
rect 2205 1124 2211 1176
rect 2237 1164 2243 1176
rect 2237 1104 2243 1156
rect 2093 957 2108 963
rect 2109 937 2140 943
rect 2093 824 2099 936
rect 2109 884 2115 937
rect 1949 724 1955 736
rect 1949 684 1955 696
rect 1709 564 1715 636
rect 1725 604 1731 656
rect 1741 644 1747 676
rect 1837 664 1843 676
rect 1981 664 1987 716
rect 2125 704 2131 836
rect 2141 704 2147 876
rect 2157 864 2163 916
rect 2173 824 2179 1080
rect 2189 1024 2195 1076
rect 2205 984 2211 996
rect 2269 983 2275 1716
rect 2301 1563 2307 2116
rect 2317 1904 2323 2156
rect 2333 1823 2339 1996
rect 2349 1983 2355 2256
rect 2461 2164 2467 2436
rect 2477 2224 2483 2256
rect 2493 2244 2499 2356
rect 2525 2323 2531 2656
rect 2557 2564 2563 2596
rect 2637 2584 2643 2716
rect 2685 2704 2691 3336
rect 2733 3204 2739 3316
rect 2717 3024 2723 3056
rect 2749 3004 2755 3636
rect 2845 3564 2851 3736
rect 2861 3484 2867 3536
rect 3021 3484 3027 4117
rect 3037 4004 3043 4076
rect 3053 4064 3059 4236
rect 3069 4143 3075 4536
rect 3149 4424 3155 4656
rect 3213 4644 3219 4696
rect 3277 4684 3283 4897
rect 3293 4684 3299 4836
rect 3309 4744 3315 4916
rect 3341 4864 3347 5237
rect 3437 5164 3443 5276
rect 3469 5263 3475 5316
rect 3492 5297 3500 5303
rect 3453 5257 3475 5263
rect 3357 5024 3363 5116
rect 3437 5084 3443 5136
rect 3453 5104 3459 5257
rect 3453 5084 3459 5096
rect 3469 5063 3475 5236
rect 3485 5124 3491 5296
rect 3565 5104 3571 5296
rect 3453 5057 3475 5063
rect 3357 4904 3363 5016
rect 3389 4984 3395 4996
rect 3437 4984 3443 5056
rect 3405 4924 3411 4936
rect 3428 4917 3443 4923
rect 3389 4704 3395 4856
rect 3389 4684 3395 4696
rect 3405 4684 3411 4916
rect 3437 4784 3443 4917
rect 3453 4844 3459 5057
rect 3469 4924 3475 4936
rect 3517 4924 3523 5036
rect 3533 4984 3539 5076
rect 3549 5024 3555 5096
rect 3581 4984 3587 5316
rect 3597 5304 3603 5457
rect 3645 5424 3651 5463
rect 3661 5457 3683 5463
rect 3613 5384 3619 5416
rect 3661 5384 3667 5457
rect 3709 5384 3715 5463
rect 3805 5457 3827 5463
rect 3597 5124 3603 5136
rect 3533 4944 3539 4976
rect 3581 4944 3587 4976
rect 3533 4924 3539 4936
rect 3453 4784 3459 4796
rect 3469 4784 3475 4896
rect 3565 4804 3571 4916
rect 3597 4904 3603 5116
rect 3629 4923 3635 5316
rect 3677 4964 3683 5316
rect 3805 5184 3811 5457
rect 5946 5414 5958 5416
rect 5931 5406 5933 5414
rect 5941 5406 5943 5414
rect 5951 5406 5953 5414
rect 5961 5406 5963 5414
rect 5971 5406 5973 5414
rect 5946 5404 5958 5406
rect 3917 5364 3923 5376
rect 4205 5364 4211 5376
rect 4317 5364 4323 5396
rect 4317 5344 4323 5356
rect 4205 5337 4220 5343
rect 3853 5326 3859 5336
rect 3885 5144 3891 5336
rect 3949 5304 3955 5316
rect 3997 5304 4003 5336
rect 4013 5124 4019 5316
rect 3629 4917 3651 4923
rect 3565 4704 3571 4756
rect 3229 4604 3235 4636
rect 3165 4526 3171 4576
rect 3101 4384 3107 4416
rect 3085 4304 3091 4356
rect 3181 4264 3187 4436
rect 3101 4224 3107 4236
rect 3181 4144 3187 4256
rect 3069 4137 3084 4143
rect 3069 4084 3075 4116
rect 3085 4104 3091 4136
rect 3085 3904 3091 3956
rect 3037 3744 3043 3896
rect 3149 3884 3155 4096
rect 3181 3904 3187 4136
rect 3197 3964 3203 4436
rect 3213 4083 3219 4276
rect 3229 4224 3235 4294
rect 3261 4184 3267 4316
rect 3309 4304 3315 4636
rect 3325 4444 3331 4636
rect 3389 4544 3395 4656
rect 3405 4604 3411 4656
rect 3357 4526 3363 4536
rect 3357 4384 3363 4496
rect 3421 4404 3427 4436
rect 3437 4404 3443 4656
rect 3501 4644 3507 4696
rect 3453 4524 3459 4616
rect 3469 4544 3475 4556
rect 3485 4544 3491 4596
rect 3517 4584 3523 4656
rect 3533 4604 3539 4636
rect 3565 4584 3571 4676
rect 3581 4624 3587 4636
rect 3645 4624 3651 4917
rect 3693 4884 3699 4916
rect 3709 4784 3715 4836
rect 3325 4304 3331 4316
rect 3405 4284 3411 4296
rect 3421 4284 3427 4396
rect 3453 4383 3459 4496
rect 3501 4384 3507 4556
rect 3444 4377 3459 4383
rect 3517 4323 3523 4496
rect 3549 4384 3555 4556
rect 3565 4544 3571 4576
rect 3565 4524 3571 4536
rect 3581 4524 3587 4596
rect 3661 4584 3667 4696
rect 3741 4684 3747 5056
rect 3773 4924 3779 5076
rect 3805 4704 3811 4796
rect 3837 4683 3843 5096
rect 3965 5063 3971 5096
rect 3981 5084 3987 5094
rect 4093 5064 4099 5336
rect 4205 5244 4211 5337
rect 4397 5324 4403 5376
rect 4557 5324 4563 5376
rect 4589 5324 4595 5356
rect 4237 5264 4243 5316
rect 4493 5303 4499 5316
rect 4292 5297 4307 5303
rect 4493 5297 4515 5303
rect 4301 5264 4307 5297
rect 3965 5057 3987 5063
rect 3860 5037 3875 5043
rect 3853 4784 3859 4836
rect 3869 4824 3875 5037
rect 3981 4984 3987 5057
rect 3965 4944 3971 4956
rect 3933 4844 3939 4916
rect 3949 4864 3955 4936
rect 3837 4677 3859 4683
rect 3693 4664 3699 4676
rect 3597 4504 3603 4516
rect 3613 4384 3619 4556
rect 3677 4544 3683 4576
rect 3693 4564 3699 4656
rect 3709 4584 3715 4616
rect 3773 4584 3779 4636
rect 3517 4317 3532 4323
rect 3341 4184 3347 4276
rect 3437 4124 3443 4296
rect 3469 4164 3475 4256
rect 3245 4104 3251 4116
rect 3213 4077 3235 4083
rect 3213 3984 3219 4036
rect 3197 3904 3203 3956
rect 3213 3884 3219 3956
rect 3149 3844 3155 3876
rect 3101 3803 3107 3836
rect 3085 3797 3107 3803
rect 3037 3724 3043 3736
rect 3037 3584 3043 3696
rect 2765 3144 2771 3336
rect 2813 3324 2819 3436
rect 2861 3364 2867 3376
rect 2829 3204 2835 3236
rect 2781 3124 2787 3196
rect 2765 3104 2771 3116
rect 2797 3084 2803 3116
rect 2861 3097 2876 3103
rect 2717 2944 2723 2976
rect 2733 2923 2739 2956
rect 2765 2924 2771 3036
rect 2781 2964 2787 3036
rect 2813 2964 2819 2976
rect 2717 2917 2739 2923
rect 2717 2784 2723 2917
rect 2829 2884 2835 3096
rect 2861 2944 2867 3097
rect 2877 2984 2883 3016
rect 2893 2964 2899 3436
rect 2938 3414 2950 3416
rect 2923 3406 2925 3414
rect 2933 3406 2935 3414
rect 2943 3406 2945 3414
rect 2953 3406 2955 3414
rect 2963 3406 2965 3414
rect 2938 3404 2950 3406
rect 2941 3344 2947 3356
rect 3053 3343 3059 3776
rect 3085 3724 3091 3797
rect 3213 3784 3219 3876
rect 3229 3844 3235 4077
rect 3325 4044 3331 4096
rect 3261 3744 3267 3836
rect 3293 3744 3299 3856
rect 3229 3726 3235 3736
rect 3181 3584 3187 3676
rect 3069 3444 3075 3480
rect 3133 3424 3139 3496
rect 3069 3364 3075 3396
rect 3261 3383 3267 3736
rect 3293 3524 3299 3736
rect 3309 3724 3315 3896
rect 3325 3664 3331 3836
rect 3341 3724 3347 3736
rect 3357 3724 3363 3736
rect 3373 3723 3379 4116
rect 3437 4084 3443 4116
rect 3437 3984 3443 4076
rect 3453 4004 3459 4136
rect 3469 4124 3475 4136
rect 3485 4124 3491 4276
rect 3501 4144 3507 4296
rect 3517 4144 3523 4216
rect 3389 3744 3395 3776
rect 3373 3717 3395 3723
rect 3389 3584 3395 3717
rect 3421 3704 3427 3836
rect 3453 3724 3459 3856
rect 3469 3704 3475 3956
rect 3453 3664 3459 3676
rect 3485 3624 3491 4116
rect 3533 3984 3539 4236
rect 3565 4064 3571 4116
rect 3565 3844 3571 3876
rect 3517 3684 3523 3776
rect 3533 3604 3539 3736
rect 3549 3704 3555 3716
rect 3277 3384 3283 3416
rect 3245 3377 3267 3383
rect 3044 3337 3059 3343
rect 2909 3184 2915 3296
rect 3053 3264 3059 3337
rect 2938 3014 2950 3016
rect 2923 3006 2925 3014
rect 2933 3006 2935 3014
rect 2943 3006 2945 3014
rect 2953 3006 2955 3014
rect 2963 3006 2965 3014
rect 2938 3004 2950 3006
rect 2909 2924 2915 2956
rect 2877 2884 2883 2916
rect 2781 2784 2787 2796
rect 2653 2684 2659 2696
rect 2717 2584 2723 2676
rect 2733 2664 2739 2736
rect 2813 2724 2819 2876
rect 2829 2724 2835 2836
rect 2941 2724 2947 2836
rect 2989 2704 2995 3116
rect 3005 3084 3011 3156
rect 3021 3104 3027 3176
rect 3053 3164 3059 3236
rect 3053 3104 3059 3136
rect 3037 3064 3043 3076
rect 3085 3024 3091 3056
rect 3021 2964 3027 2996
rect 3101 2964 3107 3236
rect 3117 3084 3123 3256
rect 3197 3143 3203 3356
rect 3245 3344 3251 3377
rect 3293 3364 3299 3476
rect 3213 3224 3219 3318
rect 3197 3137 3219 3143
rect 3213 3084 3219 3137
rect 3245 3084 3251 3336
rect 3309 3324 3315 3496
rect 3325 3324 3331 3476
rect 3421 3464 3427 3516
rect 3437 3504 3443 3596
rect 3453 3463 3459 3516
rect 3565 3504 3571 3836
rect 3581 3804 3587 4296
rect 3613 4144 3619 4296
rect 3629 4204 3635 4336
rect 3645 4324 3651 4536
rect 3757 4524 3763 4536
rect 3693 4344 3699 4516
rect 3709 4304 3715 4496
rect 3725 4304 3731 4456
rect 3757 4384 3763 4496
rect 3789 4404 3795 4556
rect 3805 4524 3811 4536
rect 3805 4423 3811 4516
rect 3837 4504 3843 4656
rect 3853 4584 3859 4677
rect 3837 4484 3843 4496
rect 3869 4464 3875 4636
rect 3805 4417 3827 4423
rect 3629 4124 3635 4196
rect 3661 4163 3667 4236
rect 3661 4157 3676 4163
rect 3693 4144 3699 4296
rect 3709 4264 3715 4276
rect 3725 4144 3731 4276
rect 3741 4184 3747 4216
rect 3677 4124 3683 4136
rect 3741 4124 3747 4176
rect 3677 4024 3683 4036
rect 3725 3964 3731 4116
rect 3741 4104 3747 4116
rect 3757 4044 3763 4236
rect 3789 4203 3795 4396
rect 3789 4197 3811 4203
rect 3661 3784 3667 3896
rect 3725 3784 3731 3896
rect 3805 3884 3811 4197
rect 3821 4184 3827 4417
rect 3885 4304 3891 4556
rect 3901 4524 3907 4536
rect 3917 4464 3923 4516
rect 3933 4484 3939 4516
rect 3949 4424 3955 4856
rect 3997 4844 4003 4936
rect 4013 4924 4019 4996
rect 4045 4984 4051 5036
rect 4093 4944 4099 5056
rect 4205 5044 4211 5236
rect 4301 5124 4307 5256
rect 4381 5124 4387 5236
rect 4442 5214 4454 5216
rect 4427 5206 4429 5214
rect 4437 5206 4439 5214
rect 4447 5206 4449 5214
rect 4457 5206 4459 5214
rect 4467 5206 4469 5214
rect 4442 5204 4454 5206
rect 4237 5084 4243 5116
rect 4141 4924 4147 4956
rect 4237 4944 4243 5076
rect 4253 5064 4259 5096
rect 4285 4984 4291 5076
rect 4301 5064 4307 5116
rect 4333 5084 4339 5096
rect 4461 5084 4467 5094
rect 4333 5044 4339 5076
rect 4365 4984 4371 5076
rect 4429 4964 4435 5036
rect 4189 4864 4195 4916
rect 4077 4704 4083 4836
rect 4077 4684 4083 4696
rect 4029 4564 4035 4676
rect 3981 4524 3987 4536
rect 4013 4504 4019 4516
rect 4061 4504 4067 4676
rect 4093 4544 4099 4556
rect 4109 4544 4115 4716
rect 4269 4704 4275 4956
rect 4445 4944 4451 4976
rect 4301 4704 4307 4936
rect 4333 4924 4339 4936
rect 4397 4924 4403 4936
rect 4317 4844 4323 4916
rect 4173 4644 4179 4696
rect 4333 4684 4339 4916
rect 4365 4704 4371 4736
rect 4349 4684 4355 4696
rect 4189 4664 4195 4676
rect 4157 4526 4163 4556
rect 3949 4384 3955 4396
rect 3965 4384 3971 4476
rect 3997 4384 4003 4456
rect 4013 4384 4019 4496
rect 4029 4364 4035 4436
rect 4237 4384 4243 4536
rect 4285 4524 4291 4576
rect 4301 4524 4307 4676
rect 4397 4643 4403 4916
rect 4493 4864 4499 5076
rect 4442 4814 4454 4816
rect 4427 4806 4429 4814
rect 4437 4806 4439 4814
rect 4447 4806 4449 4814
rect 4457 4806 4459 4814
rect 4467 4806 4469 4814
rect 4442 4804 4454 4806
rect 4493 4724 4499 4856
rect 4509 4784 4515 5297
rect 4541 5184 4547 5236
rect 4573 5164 4579 5316
rect 4621 5264 4627 5316
rect 4669 5264 4675 5336
rect 4701 5324 4707 5376
rect 5293 5344 5299 5356
rect 4797 5324 4803 5336
rect 4557 4983 4563 5056
rect 4573 5023 4579 5156
rect 4621 5104 4627 5116
rect 4573 5017 4595 5023
rect 4541 4977 4563 4983
rect 4541 4904 4547 4977
rect 4573 4964 4579 4996
rect 4589 4864 4595 5017
rect 4605 4944 4611 4996
rect 4621 4944 4627 5036
rect 4605 4904 4611 4916
rect 4525 4744 4531 4816
rect 4621 4784 4627 4916
rect 4605 4777 4620 4783
rect 4493 4664 4499 4716
rect 4397 4637 4419 4643
rect 4333 4564 4339 4636
rect 4397 4564 4403 4576
rect 4413 4524 4419 4637
rect 3837 4184 3843 4296
rect 3965 4144 3971 4256
rect 3981 4184 3987 4256
rect 3821 4084 3827 4116
rect 3949 3984 3955 4136
rect 3997 3984 4003 4116
rect 4013 4084 4019 4256
rect 4029 4204 4035 4236
rect 4189 4223 4195 4296
rect 4173 4217 4195 4223
rect 4093 4144 4099 4216
rect 4173 4184 4179 4217
rect 4237 4184 4243 4276
rect 3821 3924 3827 3976
rect 3988 3917 4003 3923
rect 3805 3864 3811 3876
rect 3741 3844 3747 3856
rect 3597 3724 3603 3776
rect 3757 3764 3763 3856
rect 3789 3784 3795 3836
rect 3837 3784 3843 3836
rect 3853 3804 3859 3876
rect 3652 3737 3683 3743
rect 3613 3717 3628 3723
rect 3597 3524 3603 3696
rect 3613 3684 3619 3717
rect 3677 3703 3683 3737
rect 3741 3724 3747 3736
rect 3773 3724 3779 3776
rect 3821 3724 3827 3756
rect 3757 3704 3763 3716
rect 3677 3697 3708 3703
rect 3597 3484 3603 3496
rect 3453 3457 3475 3463
rect 3389 3384 3395 3456
rect 3453 3444 3459 3457
rect 3389 3324 3395 3376
rect 3309 3204 3315 3316
rect 3469 3304 3475 3457
rect 3485 3384 3491 3456
rect 3405 3284 3411 3296
rect 3133 2964 3139 2976
rect 3069 2924 3075 2956
rect 3149 2904 3155 3036
rect 3213 3004 3219 3076
rect 3293 3044 3299 3096
rect 3277 2944 3283 2956
rect 3229 2904 3235 2936
rect 3309 2924 3315 3196
rect 3245 2884 3251 2916
rect 3053 2824 3059 2876
rect 3261 2864 3267 2916
rect 3341 2904 3347 3136
rect 3373 2984 3379 3276
rect 3437 3264 3443 3276
rect 3421 3184 3427 3216
rect 3405 3104 3411 3136
rect 3453 3084 3459 3156
rect 3469 3144 3475 3296
rect 3501 3144 3507 3416
rect 3517 3344 3523 3476
rect 3613 3384 3619 3636
rect 3677 3484 3683 3496
rect 3725 3484 3731 3556
rect 3741 3504 3747 3656
rect 3757 3584 3763 3696
rect 3645 3444 3651 3476
rect 3741 3464 3747 3476
rect 3789 3463 3795 3496
rect 3805 3484 3811 3716
rect 3837 3504 3843 3756
rect 3869 3724 3875 3876
rect 3885 3844 3891 3896
rect 3933 3864 3939 3876
rect 3901 3744 3907 3796
rect 3997 3784 4003 3917
rect 3853 3704 3859 3716
rect 3869 3524 3875 3616
rect 3837 3464 3843 3496
rect 3853 3464 3859 3516
rect 3789 3457 3811 3463
rect 3549 3344 3555 3356
rect 3677 3344 3683 3396
rect 3741 3344 3747 3436
rect 3549 3284 3555 3336
rect 3661 3304 3667 3316
rect 3613 3264 3619 3296
rect 3533 3163 3539 3236
rect 3629 3184 3635 3196
rect 3533 3157 3555 3163
rect 3533 3124 3539 3136
rect 3549 3124 3555 3157
rect 3709 3124 3715 3136
rect 3405 2964 3411 3076
rect 3421 2984 3427 3056
rect 3437 2984 3443 3056
rect 2829 2584 2835 2656
rect 2509 2317 2531 2323
rect 2509 2184 2515 2317
rect 2541 2304 2547 2316
rect 2557 2284 2563 2536
rect 2573 2284 2579 2376
rect 2669 2324 2675 2536
rect 2685 2283 2691 2536
rect 2701 2284 2707 2436
rect 2676 2277 2691 2283
rect 2525 2164 2531 2216
rect 2541 2184 2547 2256
rect 2605 2224 2611 2236
rect 2621 2184 2627 2216
rect 2669 2164 2675 2276
rect 2701 2264 2707 2276
rect 2685 2164 2691 2176
rect 2717 2164 2723 2516
rect 2749 2324 2755 2356
rect 2749 2184 2755 2276
rect 2365 2124 2371 2136
rect 2372 2057 2403 2063
rect 2397 2044 2403 2057
rect 2349 1977 2371 1983
rect 2317 1817 2339 1823
rect 2317 1744 2323 1817
rect 2349 1763 2355 1956
rect 2365 1924 2371 1977
rect 2381 1904 2387 2036
rect 2413 1923 2419 2056
rect 2429 1924 2435 2096
rect 2397 1917 2419 1923
rect 2397 1844 2403 1917
rect 2413 1784 2419 1856
rect 2340 1757 2355 1763
rect 2333 1723 2339 1736
rect 2317 1717 2339 1723
rect 2349 1723 2355 1736
rect 2349 1717 2364 1723
rect 2317 1584 2323 1717
rect 2349 1584 2355 1656
rect 2365 1644 2371 1716
rect 2301 1557 2323 1563
rect 2317 1464 2323 1557
rect 2445 1524 2451 2056
rect 2509 2024 2515 2096
rect 2461 1944 2467 2016
rect 2541 1963 2547 2156
rect 2669 2124 2675 2136
rect 2557 2104 2563 2116
rect 2541 1957 2563 1963
rect 2461 1784 2467 1876
rect 2477 1784 2483 1916
rect 2493 1904 2499 1916
rect 2541 1823 2547 1916
rect 2557 1904 2563 1957
rect 2525 1817 2547 1823
rect 2525 1784 2531 1817
rect 2461 1704 2467 1716
rect 2509 1684 2515 1756
rect 2525 1737 2540 1743
rect 2525 1664 2531 1737
rect 2541 1704 2547 1716
rect 2557 1584 2563 1876
rect 2605 1844 2611 1856
rect 2573 1724 2579 1736
rect 2621 1584 2627 1736
rect 2621 1544 2627 1576
rect 2301 1384 2307 1456
rect 2317 1363 2323 1456
rect 2333 1444 2339 1456
rect 2349 1364 2355 1516
rect 2365 1384 2371 1456
rect 2301 1357 2323 1363
rect 2301 1184 2307 1357
rect 2333 1304 2339 1336
rect 2381 1324 2387 1496
rect 2413 1384 2419 1496
rect 2429 1484 2435 1496
rect 2461 1404 2467 1496
rect 2477 1484 2483 1496
rect 2525 1483 2531 1496
rect 2493 1404 2499 1480
rect 2525 1477 2540 1483
rect 2557 1464 2563 1496
rect 2397 1264 2403 1316
rect 2445 1264 2451 1316
rect 2285 1004 2291 1096
rect 2301 1084 2307 1176
rect 2333 1064 2339 1096
rect 2269 977 2284 983
rect 2253 924 2259 976
rect 2269 864 2275 936
rect 2301 763 2307 916
rect 2333 824 2339 956
rect 2317 784 2323 816
rect 2301 757 2323 763
rect 2237 704 2243 716
rect 2253 684 2259 756
rect 2269 683 2275 696
rect 2269 677 2291 683
rect 1725 564 1731 596
rect 1741 564 1747 636
rect 1837 604 1843 656
rect 1789 584 1795 596
rect 1773 544 1779 556
rect 1869 544 1875 596
rect 1949 564 1955 596
rect 1549 304 1555 376
rect 1581 304 1587 496
rect 1645 384 1651 476
rect 1757 384 1763 456
rect 1837 324 1843 336
rect 1853 324 1859 436
rect 1869 384 1875 536
rect 1965 524 1971 636
rect 1981 544 1987 656
rect 1997 564 2003 676
rect 2093 664 2099 676
rect 2109 563 2115 636
rect 2100 557 2115 563
rect 2029 544 2035 556
rect 2141 544 2147 576
rect 2189 564 2195 636
rect 2205 584 2211 616
rect 2221 564 2227 676
rect 2157 524 2163 556
rect 1604 317 1619 323
rect 1597 284 1603 296
rect 1613 284 1619 317
rect 1917 304 1923 436
rect 2157 384 2163 496
rect 1709 284 1715 296
rect 1533 244 1539 276
rect 1533 144 1539 176
rect 909 124 915 136
rect 1117 124 1123 136
rect 381 103 387 116
rect 493 104 499 116
rect 1133 104 1139 136
rect 1549 104 1555 156
rect 1597 144 1603 256
rect 1613 204 1619 236
rect 1645 184 1651 236
rect 1661 224 1667 256
rect 372 97 387 103
rect 445 84 451 96
rect 461 84 467 96
rect 1277 84 1283 96
rect 1661 84 1667 196
rect 1709 164 1715 216
rect 1757 164 1763 256
rect 1773 184 1779 276
rect 1789 163 1795 296
rect 1805 184 1811 296
rect 1837 184 1843 296
rect 1869 204 1875 276
rect 1917 244 1923 296
rect 1965 284 1971 376
rect 1805 164 1811 176
rect 1773 157 1795 163
rect 1693 104 1699 136
rect 1773 104 1779 157
rect 1885 144 1891 216
rect 1965 164 1971 256
rect 1981 244 1987 256
rect 1997 204 2003 236
rect 1965 144 1971 156
rect 1997 144 2003 176
rect 2013 164 2019 296
rect 2029 284 2035 356
rect 2093 337 2147 343
rect 2093 324 2099 337
rect 2141 324 2147 337
rect 2125 284 2131 316
rect 2189 284 2195 536
rect 2221 503 2227 516
rect 2221 497 2243 503
rect 2237 384 2243 497
rect 2205 304 2211 376
rect 2029 184 2035 256
rect 2141 244 2147 256
rect 2077 164 2083 196
rect 2157 144 2163 256
rect 2189 164 2195 236
rect 2237 204 2243 336
rect 2253 304 2259 476
rect 2269 384 2275 656
rect 2285 604 2291 677
rect 2301 644 2307 736
rect 2301 524 2307 636
rect 2317 524 2323 757
rect 2349 703 2355 996
rect 2365 984 2371 1256
rect 2397 1184 2403 1196
rect 2461 1184 2467 1396
rect 2525 1384 2531 1436
rect 2573 1364 2579 1496
rect 2589 1484 2595 1496
rect 2605 1384 2611 1396
rect 2637 1384 2643 2096
rect 2733 2064 2739 2096
rect 2669 1984 2675 2016
rect 2685 1804 2691 1864
rect 2653 1764 2659 1796
rect 2733 1784 2739 1876
rect 2749 1764 2755 2156
rect 2765 2144 2771 2476
rect 2781 2384 2787 2536
rect 2813 2504 2819 2556
rect 2781 2344 2787 2376
rect 2797 2323 2803 2456
rect 2845 2384 2851 2496
rect 2788 2317 2803 2323
rect 2861 2304 2867 2696
rect 2938 2614 2950 2616
rect 2923 2606 2925 2614
rect 2933 2606 2935 2614
rect 2943 2606 2945 2614
rect 2953 2606 2955 2614
rect 2963 2606 2965 2614
rect 2938 2604 2950 2606
rect 2973 2324 2979 2436
rect 2989 2404 2995 2556
rect 3069 2543 3075 2836
rect 3101 2684 3107 2696
rect 3085 2624 3091 2676
rect 3117 2604 3123 2836
rect 3149 2784 3155 2836
rect 3117 2564 3123 2576
rect 3133 2564 3139 2776
rect 3197 2704 3203 2836
rect 3069 2537 3091 2543
rect 3085 2524 3091 2537
rect 3101 2524 3107 2536
rect 3005 2364 3011 2436
rect 3053 2324 3059 2356
rect 2909 2244 2915 2276
rect 2845 2184 2851 2236
rect 2938 2214 2950 2216
rect 2923 2206 2925 2214
rect 2933 2206 2935 2214
rect 2943 2206 2945 2214
rect 2953 2206 2955 2214
rect 2963 2206 2965 2214
rect 2938 2204 2950 2206
rect 3037 2184 3043 2276
rect 3053 2163 3059 2236
rect 3069 2184 3075 2516
rect 3149 2344 3155 2596
rect 3197 2544 3203 2616
rect 3117 2324 3123 2336
rect 3165 2324 3171 2436
rect 3197 2384 3203 2396
rect 3229 2324 3235 2776
rect 3245 2684 3251 2716
rect 3261 2524 3267 2676
rect 3277 2664 3283 2776
rect 3341 2724 3347 2896
rect 3357 2864 3363 2916
rect 3373 2744 3379 2756
rect 3405 2704 3411 2956
rect 3421 2784 3427 2976
rect 3469 2964 3475 3096
rect 3501 2984 3507 3036
rect 3485 2964 3491 2976
rect 3453 2924 3459 2956
rect 3469 2944 3475 2956
rect 3517 2944 3523 3016
rect 3533 2943 3539 3116
rect 3565 3097 3580 3103
rect 3533 2937 3555 2943
rect 3469 2904 3475 2936
rect 3533 2904 3539 2916
rect 3549 2904 3555 2937
rect 3565 2924 3571 3097
rect 3597 3064 3603 3076
rect 3613 2944 3619 3116
rect 3629 3084 3635 3096
rect 3645 3004 3651 3076
rect 3661 2944 3667 2956
rect 3677 2944 3683 3076
rect 3709 3044 3715 3116
rect 3725 3104 3731 3276
rect 3805 3184 3811 3457
rect 3869 3304 3875 3436
rect 3885 3284 3891 3716
rect 3901 3484 3907 3736
rect 3917 3504 3923 3696
rect 3949 3664 3955 3676
rect 3933 3484 3939 3556
rect 3981 3504 3987 3576
rect 3997 3564 4003 3736
rect 4013 3544 4019 4036
rect 4061 3884 4067 4136
rect 4093 3984 4099 4136
rect 4109 4124 4115 4156
rect 4189 4144 4195 4156
rect 4141 4104 4147 4116
rect 4205 4104 4211 4116
rect 4061 3764 4067 3876
rect 4077 3864 4083 3896
rect 4029 3724 4035 3736
rect 4045 3704 4051 3716
rect 3997 3524 4003 3536
rect 4045 3504 4051 3696
rect 4077 3684 4083 3856
rect 4125 3804 4131 4076
rect 4189 3924 4195 3976
rect 4141 3784 4147 3896
rect 4221 3784 4227 3996
rect 4269 3924 4275 4516
rect 4333 4284 4339 4516
rect 4442 4414 4454 4416
rect 4427 4406 4429 4414
rect 4437 4406 4439 4414
rect 4447 4406 4449 4414
rect 4457 4406 4459 4414
rect 4467 4406 4469 4414
rect 4442 4404 4454 4406
rect 4493 4284 4499 4656
rect 4589 4544 4595 4656
rect 4557 4524 4563 4536
rect 4605 4524 4611 4777
rect 4637 4744 4643 5216
rect 4685 5144 4691 5316
rect 4660 5117 4707 5123
rect 4701 5104 4707 5117
rect 4749 5104 4755 5116
rect 4797 5104 4803 5176
rect 4685 5083 4691 5096
rect 4685 5077 4707 5083
rect 4653 4963 4659 5076
rect 4669 4984 4675 5076
rect 4701 5044 4707 5077
rect 4653 4957 4675 4963
rect 4669 4904 4675 4957
rect 4685 4944 4691 5036
rect 4717 5024 4723 5036
rect 4733 4984 4739 5016
rect 4749 4924 4755 4996
rect 4765 4944 4771 4956
rect 4653 4824 4659 4896
rect 4669 4824 4675 4896
rect 4685 4864 4691 4916
rect 4733 4864 4739 4896
rect 4781 4863 4787 5076
rect 4797 5004 4803 5036
rect 4813 5004 4819 5336
rect 4829 4924 4835 5316
rect 4909 5204 4915 5316
rect 4957 5304 4963 5316
rect 4989 5244 4995 5336
rect 5053 5324 5059 5336
rect 5005 5224 5011 5316
rect 5053 5224 5059 5296
rect 5085 5284 5091 5336
rect 5341 5324 5347 5356
rect 5357 5304 5363 5336
rect 5565 5326 5571 5356
rect 5629 5344 5635 5376
rect 5021 5184 5027 5196
rect 5085 5184 5091 5276
rect 4893 5104 4899 5116
rect 5117 5104 5123 5156
rect 5149 5104 5155 5116
rect 4868 5097 4883 5103
rect 4877 5083 4883 5097
rect 5229 5103 5235 5116
rect 5229 5097 5244 5103
rect 4877 5077 4892 5083
rect 4845 5024 4851 5076
rect 4861 5064 4867 5076
rect 4909 5064 4915 5076
rect 4957 5004 4963 5096
rect 4861 4944 4867 4996
rect 4989 4984 4995 5056
rect 5053 5024 5059 5096
rect 5069 5063 5075 5076
rect 5069 5057 5091 5063
rect 5021 4964 5027 4976
rect 5069 4964 5075 5036
rect 4772 4857 4787 4863
rect 4637 4704 4643 4736
rect 4653 4704 4659 4716
rect 4669 4603 4675 4816
rect 4685 4664 4691 4856
rect 4701 4724 4707 4736
rect 4733 4684 4739 4756
rect 4653 4597 4675 4603
rect 4653 4544 4659 4597
rect 4733 4584 4739 4656
rect 4749 4644 4755 4656
rect 4765 4644 4771 4856
rect 4813 4764 4819 4916
rect 4781 4564 4787 4656
rect 4637 4524 4643 4536
rect 4717 4524 4723 4536
rect 4813 4524 4819 4736
rect 4285 3984 4291 3996
rect 4317 3944 4323 4256
rect 4349 4144 4355 4276
rect 4509 4184 4515 4296
rect 4237 3804 4243 3876
rect 4253 3784 4259 3916
rect 4269 3823 4275 3836
rect 4269 3817 4291 3823
rect 4093 3724 4099 3776
rect 4221 3764 4227 3776
rect 4109 3704 4115 3756
rect 4125 3684 4131 3716
rect 4093 3544 4099 3636
rect 4077 3524 4083 3536
rect 4109 3504 4115 3676
rect 4141 3584 4147 3676
rect 3917 3477 3932 3483
rect 3917 3343 3923 3477
rect 3933 3384 3939 3396
rect 3917 3337 3932 3343
rect 3773 3124 3779 3156
rect 3789 3104 3795 3116
rect 3693 2984 3699 3016
rect 3677 2924 3683 2936
rect 3613 2904 3619 2916
rect 3629 2904 3635 2916
rect 3325 2684 3331 2696
rect 3309 2663 3315 2676
rect 3309 2657 3331 2663
rect 3277 2564 3283 2656
rect 3325 2584 3331 2657
rect 3405 2644 3411 2696
rect 3293 2504 3299 2516
rect 3373 2444 3379 2536
rect 3373 2324 3379 2436
rect 3053 2157 3075 2163
rect 2765 2064 2771 2136
rect 2781 1964 2787 2136
rect 2845 2024 2851 2076
rect 2788 1957 2803 1963
rect 2765 1764 2771 1896
rect 2797 1744 2803 1957
rect 2813 1944 2819 1956
rect 2861 1924 2867 2076
rect 2877 2004 2883 2136
rect 3053 2004 3059 2136
rect 3069 2084 3075 2157
rect 2877 1937 2915 1943
rect 2813 1864 2819 1916
rect 2877 1903 2883 1937
rect 2909 1923 2915 1937
rect 2909 1917 2924 1923
rect 2868 1897 2883 1903
rect 2829 1784 2835 1896
rect 3053 1863 3059 1916
rect 3085 1904 3091 2296
rect 3101 1884 3107 2276
rect 3373 2244 3379 2296
rect 3117 2164 3123 2236
rect 3229 2224 3235 2236
rect 3229 2144 3235 2216
rect 3213 2124 3219 2136
rect 3261 2124 3267 2236
rect 3293 2117 3308 2123
rect 3133 1864 3139 1936
rect 3037 1857 3059 1863
rect 2845 1824 2851 1856
rect 2717 1724 2723 1736
rect 2781 1724 2787 1736
rect 2701 1624 2707 1716
rect 2653 1504 2659 1556
rect 2717 1504 2723 1716
rect 2765 1624 2771 1716
rect 2797 1624 2803 1716
rect 2829 1584 2835 1756
rect 2845 1744 2851 1796
rect 2877 1784 2883 1856
rect 3037 1844 3043 1857
rect 2938 1814 2950 1816
rect 2923 1806 2925 1814
rect 2933 1806 2935 1814
rect 2943 1806 2945 1814
rect 2953 1806 2955 1814
rect 2963 1806 2965 1814
rect 2938 1804 2950 1806
rect 2941 1744 2947 1776
rect 2845 1724 2851 1736
rect 2813 1524 2819 1536
rect 2701 1484 2707 1496
rect 2813 1484 2819 1516
rect 2845 1497 2860 1503
rect 2557 1344 2563 1356
rect 2573 1344 2579 1356
rect 2669 1344 2675 1456
rect 2717 1403 2723 1436
rect 2717 1397 2739 1403
rect 2701 1344 2707 1396
rect 2733 1344 2739 1397
rect 2749 1384 2755 1416
rect 2765 1344 2771 1456
rect 2493 1304 2499 1316
rect 2461 1104 2467 1116
rect 2429 1044 2435 1076
rect 2461 984 2467 1076
rect 2493 1024 2499 1296
rect 2509 1184 2515 1196
rect 2525 1184 2531 1296
rect 2557 1283 2563 1336
rect 2605 1304 2611 1336
rect 2541 1277 2563 1283
rect 2541 1083 2547 1277
rect 2541 1077 2563 1083
rect 2493 984 2499 1016
rect 2381 924 2387 956
rect 2429 864 2435 956
rect 2413 784 2419 856
rect 2445 764 2451 916
rect 2477 864 2483 956
rect 2493 804 2499 836
rect 2349 697 2364 703
rect 2269 283 2275 356
rect 2260 277 2275 283
rect 1853 124 1859 136
rect 2141 124 2147 136
rect 2237 124 2243 196
rect 2253 123 2259 156
rect 2285 144 2291 516
rect 2301 304 2307 476
rect 2317 384 2323 516
rect 2333 423 2339 656
rect 2349 484 2355 697
rect 2381 664 2387 736
rect 2477 724 2483 756
rect 2493 724 2499 736
rect 2413 704 2419 716
rect 2413 603 2419 656
rect 2397 597 2419 603
rect 2372 557 2387 563
rect 2365 524 2371 536
rect 2333 417 2348 423
rect 2349 304 2355 416
rect 2381 344 2387 557
rect 2397 544 2403 597
rect 2445 584 2451 656
rect 2461 584 2467 716
rect 2477 564 2483 696
rect 2509 584 2515 1056
rect 2541 944 2547 1016
rect 2541 924 2547 936
rect 2525 664 2531 796
rect 2557 704 2563 1077
rect 2589 924 2595 1256
rect 2621 1204 2627 1336
rect 2669 1324 2675 1336
rect 2797 1324 2803 1436
rect 2765 1264 2771 1316
rect 2845 1244 2851 1497
rect 2877 1324 2883 1676
rect 2893 1344 2899 1716
rect 2957 1564 2963 1636
rect 2989 1604 2995 1836
rect 2957 1544 2963 1556
rect 3037 1504 3043 1796
rect 3053 1544 3059 1836
rect 3149 1704 3155 1836
rect 3069 1523 3075 1636
rect 3053 1517 3075 1523
rect 2938 1414 2950 1416
rect 2923 1406 2925 1414
rect 2933 1406 2935 1414
rect 2943 1406 2945 1414
rect 2953 1406 2955 1414
rect 2963 1406 2965 1414
rect 2938 1404 2950 1406
rect 3005 1384 3011 1436
rect 2621 1184 2627 1196
rect 2829 1104 2835 1236
rect 2861 1124 2867 1296
rect 2893 1124 2899 1336
rect 2909 1324 2915 1336
rect 2909 1264 2915 1316
rect 2909 1104 2915 1256
rect 3021 1224 3027 1236
rect 3053 1164 3059 1517
rect 3101 1484 3107 1676
rect 3165 1624 3171 2116
rect 3213 1924 3219 2036
rect 3277 2004 3283 2096
rect 3101 1364 3107 1476
rect 3133 1444 3139 1456
rect 3181 1444 3187 1856
rect 3229 1744 3235 1976
rect 3277 1924 3283 1956
rect 3277 1724 3283 1736
rect 3245 1524 3251 1616
rect 3293 1504 3299 2117
rect 3341 1984 3347 2236
rect 3389 2024 3395 2416
rect 3405 2204 3411 2636
rect 3437 2504 3443 2516
rect 3437 2443 3443 2496
rect 3421 2437 3443 2443
rect 3421 2284 3427 2437
rect 3453 2424 3459 2676
rect 3469 2424 3475 2696
rect 3485 2684 3491 2876
rect 3565 2864 3571 2896
rect 3581 2884 3587 2896
rect 3597 2764 3603 2796
rect 3645 2784 3651 2916
rect 3549 2724 3555 2756
rect 3485 2444 3491 2676
rect 3549 2664 3555 2716
rect 3581 2704 3587 2736
rect 3597 2724 3603 2756
rect 3677 2724 3683 2756
rect 3581 2564 3587 2696
rect 3597 2684 3603 2696
rect 3709 2683 3715 2996
rect 3725 2923 3731 3056
rect 3741 2944 3747 3076
rect 3773 3004 3779 3076
rect 3789 3064 3795 3096
rect 3853 3064 3859 3136
rect 3789 2984 3795 3036
rect 3837 3024 3843 3036
rect 3837 2964 3843 3016
rect 3901 3004 3907 3056
rect 3725 2917 3740 2923
rect 3741 2904 3747 2916
rect 3757 2784 3763 2936
rect 3773 2804 3779 2956
rect 3789 2944 3795 2956
rect 3901 2924 3907 2996
rect 3933 2944 3939 3336
rect 3949 3324 3955 3456
rect 3965 3344 3971 3356
rect 3981 3324 3987 3496
rect 3997 3384 4003 3476
rect 4013 3384 4019 3436
rect 4045 3344 4051 3476
rect 3949 3104 3955 3316
rect 3981 3124 3987 3316
rect 4029 3204 4035 3316
rect 4077 3303 4083 3436
rect 4093 3304 4099 3316
rect 4068 3297 4083 3303
rect 4061 3184 4067 3276
rect 4125 3104 4131 3496
rect 4157 3484 4163 3736
rect 4237 3724 4243 3756
rect 4269 3723 4275 3796
rect 4285 3724 4291 3817
rect 4301 3744 4307 3776
rect 4317 3724 4323 3856
rect 4349 3804 4355 4136
rect 4477 4124 4483 4156
rect 4493 4124 4499 4136
rect 4442 4014 4454 4016
rect 4427 4006 4429 4014
rect 4437 4006 4439 4014
rect 4447 4006 4449 4014
rect 4457 4006 4459 4014
rect 4467 4006 4469 4014
rect 4442 4004 4454 4006
rect 4413 3804 4419 3856
rect 4445 3823 4451 3896
rect 4429 3817 4451 3823
rect 4429 3784 4435 3817
rect 4253 3717 4275 3723
rect 4205 3524 4211 3636
rect 4221 3524 4227 3636
rect 4157 3363 4163 3476
rect 4157 3357 4172 3363
rect 4205 3344 4211 3516
rect 4221 3324 4227 3496
rect 4253 3484 4259 3717
rect 4301 3704 4307 3716
rect 4301 3623 4307 3696
rect 4301 3617 4323 3623
rect 4237 3364 4243 3436
rect 4253 3344 4259 3476
rect 4301 3384 4307 3596
rect 4285 3304 4291 3376
rect 4269 3184 4275 3236
rect 4317 3184 4323 3617
rect 4365 3384 4371 3736
rect 4381 3704 4387 3716
rect 4397 3684 4403 3716
rect 4445 3664 4451 3756
rect 4477 3704 4483 3836
rect 4333 3284 4339 3316
rect 4365 3304 4371 3356
rect 4381 3184 4387 3656
rect 4442 3614 4454 3616
rect 4427 3606 4429 3614
rect 4437 3606 4439 3614
rect 4447 3606 4449 3614
rect 4457 3606 4459 3614
rect 4467 3606 4469 3614
rect 4442 3604 4454 3606
rect 4397 3484 4403 3496
rect 4413 3344 4419 3556
rect 4477 3504 4483 3576
rect 4397 3304 4403 3316
rect 4477 3304 4483 3496
rect 4493 3484 4499 4116
rect 4509 3964 4515 4016
rect 4525 4004 4531 4436
rect 4573 4164 4579 4236
rect 4589 4223 4595 4516
rect 4605 4303 4611 4516
rect 4669 4384 4675 4516
rect 4701 4504 4707 4516
rect 4765 4484 4771 4516
rect 4813 4504 4819 4516
rect 4829 4484 4835 4916
rect 4861 4723 4867 4936
rect 4909 4924 4915 4936
rect 5069 4924 5075 4936
rect 5037 4864 5043 4916
rect 5085 4864 5091 5057
rect 5133 5044 5139 5076
rect 5117 4963 5123 4996
rect 5101 4957 5123 4963
rect 4852 4717 4867 4723
rect 4845 4684 4851 4716
rect 4877 4702 4883 4716
rect 5005 4664 5011 4716
rect 5101 4704 5107 4957
rect 5117 4924 5123 4936
rect 5133 4924 5139 4936
rect 5037 4684 5043 4696
rect 5117 4684 5123 4856
rect 5149 4744 5155 5096
rect 5213 5084 5219 5096
rect 5181 4984 5187 5056
rect 5197 5044 5203 5076
rect 5309 5064 5315 5096
rect 5325 5084 5331 5116
rect 5165 4944 5171 4956
rect 5165 4764 5171 4916
rect 5213 4904 5219 4916
rect 5165 4737 5212 4743
rect 5053 4643 5059 4676
rect 5117 4664 5123 4676
rect 5053 4637 5075 4643
rect 4845 4524 4851 4556
rect 4765 4384 4771 4396
rect 4813 4324 4819 4476
rect 4877 4384 4883 4576
rect 4925 4544 4931 4636
rect 4941 4524 4947 4576
rect 4957 4544 4963 4556
rect 4813 4304 4819 4316
rect 4893 4304 4899 4496
rect 4909 4484 4915 4516
rect 4605 4297 4620 4303
rect 4637 4244 4643 4296
rect 4589 4217 4611 4223
rect 4589 4184 4595 4196
rect 4605 4124 4611 4217
rect 4653 4124 4659 4276
rect 4733 4204 4739 4296
rect 4781 4244 4787 4296
rect 4845 4284 4851 4296
rect 4717 4126 4723 4176
rect 4781 4144 4787 4196
rect 4877 4144 4883 4156
rect 4893 4124 4899 4156
rect 4861 4104 4867 4116
rect 4557 3704 4563 3716
rect 4573 3564 4579 3736
rect 4589 3704 4595 3716
rect 4605 3684 4611 3796
rect 4653 3744 4659 3976
rect 4733 3904 4739 3976
rect 4669 3744 4675 3856
rect 4701 3823 4707 3896
rect 4781 3884 4787 4096
rect 4765 3844 4771 3856
rect 4685 3817 4707 3823
rect 4685 3784 4691 3817
rect 4749 3804 4755 3836
rect 4797 3804 4803 3896
rect 4701 3764 4707 3796
rect 4493 3424 4499 3476
rect 4605 3464 4611 3676
rect 4509 3344 4515 3436
rect 4525 3404 4531 3456
rect 4541 3324 4547 3416
rect 4557 3384 4563 3396
rect 4573 3364 4579 3376
rect 4605 3344 4611 3456
rect 4621 3424 4627 3716
rect 4653 3584 4659 3716
rect 4653 3504 4659 3576
rect 4669 3502 4675 3536
rect 4701 3484 4707 3736
rect 4733 3684 4739 3736
rect 4781 3724 4787 3736
rect 4813 3624 4819 4096
rect 4861 3904 4867 4076
rect 4845 3864 4851 3896
rect 4861 3884 4867 3896
rect 4877 3644 4883 4116
rect 4909 4084 4915 4476
rect 4925 4164 4931 4176
rect 4941 4084 4947 4256
rect 4973 4164 4979 4616
rect 4989 4384 4995 4516
rect 5005 4464 5011 4496
rect 5021 4404 5027 4556
rect 5037 4484 5043 4516
rect 4989 4284 4995 4336
rect 5037 4304 5043 4476
rect 5053 4404 5059 4516
rect 5069 4444 5075 4637
rect 5133 4564 5139 4696
rect 5165 4683 5171 4737
rect 5181 4704 5187 4716
rect 5213 4704 5219 4716
rect 5165 4677 5180 4683
rect 5197 4604 5203 4676
rect 5229 4564 5235 4916
rect 5261 4784 5267 5056
rect 5325 4903 5331 5076
rect 5341 5064 5347 5196
rect 5373 5184 5379 5276
rect 5405 5164 5411 5316
rect 5357 5104 5363 5136
rect 5373 5044 5379 5136
rect 5405 5064 5411 5096
rect 5453 4963 5459 5236
rect 5469 5084 5475 5096
rect 5485 5084 5491 5176
rect 5501 5104 5507 5156
rect 5517 4964 5523 5316
rect 5629 5284 5635 5336
rect 5661 5304 5667 5316
rect 5661 5224 5667 5296
rect 5725 5224 5731 5336
rect 5757 5324 5763 5376
rect 5805 5324 5811 5356
rect 5853 5324 5859 5376
rect 5997 5364 6003 5376
rect 5901 5324 5907 5356
rect 6125 5326 6131 5336
rect 5821 5304 5827 5316
rect 5581 5104 5587 5176
rect 5437 4957 5459 4963
rect 5357 4924 5363 4956
rect 5437 4944 5443 4957
rect 5517 4944 5523 4956
rect 5309 4897 5331 4903
rect 5309 4824 5315 4897
rect 5309 4784 5315 4816
rect 5421 4764 5427 4936
rect 5245 4664 5251 4716
rect 5293 4644 5299 4696
rect 5309 4563 5315 4636
rect 5325 4584 5331 4656
rect 5293 4557 5315 4563
rect 5085 4524 5091 4536
rect 5149 4524 5155 4536
rect 5245 4524 5251 4536
rect 5069 4304 5075 4376
rect 5085 4323 5091 4436
rect 5149 4344 5155 4516
rect 5229 4484 5235 4516
rect 5085 4317 5107 4323
rect 5005 4204 5011 4296
rect 5021 4264 5027 4296
rect 4973 4144 4979 4156
rect 4957 4104 4963 4116
rect 5053 4104 5059 4118
rect 4909 3984 4915 4056
rect 4893 3824 4899 3896
rect 4909 3763 4915 3916
rect 4941 3904 4947 3936
rect 5053 3923 5059 3936
rect 5037 3917 5059 3923
rect 4989 3904 4995 3916
rect 5021 3883 5027 3916
rect 5037 3904 5043 3917
rect 5085 3904 5091 4296
rect 5101 4284 5107 4317
rect 5165 4303 5171 4436
rect 5213 4384 5219 4416
rect 5156 4297 5171 4303
rect 5117 4284 5123 4296
rect 5133 4264 5139 4276
rect 5181 4243 5187 4276
rect 5197 4264 5203 4296
rect 5181 4237 5203 4243
rect 5021 3877 5036 3883
rect 4973 3864 4979 3876
rect 4957 3843 4963 3856
rect 4957 3837 4988 3843
rect 4973 3784 4979 3816
rect 4893 3757 4915 3763
rect 4765 3524 4771 3616
rect 4813 3504 4819 3516
rect 4829 3484 4835 3496
rect 4442 3214 4454 3216
rect 4427 3206 4429 3214
rect 4437 3206 4439 3214
rect 4447 3206 4449 3214
rect 4457 3206 4459 3214
rect 4467 3206 4469 3214
rect 4442 3204 4454 3206
rect 4205 3144 4211 3176
rect 4221 3143 4227 3156
rect 4221 3137 4268 3143
rect 4237 3104 4243 3116
rect 4285 3104 4291 3116
rect 3981 3044 3987 3076
rect 4077 3024 4083 3056
rect 3965 2924 3971 2956
rect 3693 2677 3715 2683
rect 3645 2604 3651 2676
rect 3661 2664 3667 2676
rect 3645 2584 3651 2596
rect 3661 2564 3667 2656
rect 3629 2544 3635 2556
rect 3597 2444 3603 2536
rect 3629 2504 3635 2516
rect 3645 2483 3651 2556
rect 3661 2524 3667 2536
rect 3629 2477 3651 2483
rect 3437 2223 3443 2294
rect 3469 2264 3475 2356
rect 3437 2217 3459 2223
rect 3453 2204 3459 2217
rect 3405 2164 3411 2176
rect 3437 2164 3443 2196
rect 3453 2064 3459 2156
rect 3501 2144 3507 2276
rect 3517 2164 3523 2436
rect 3629 2384 3635 2477
rect 3693 2423 3699 2677
rect 3725 2664 3731 2696
rect 3709 2644 3715 2656
rect 3741 2643 3747 2756
rect 3805 2744 3811 2916
rect 3917 2897 3948 2903
rect 3885 2884 3891 2896
rect 3725 2637 3747 2643
rect 3725 2544 3731 2637
rect 3821 2623 3827 2876
rect 3837 2702 3843 2736
rect 3821 2617 3843 2623
rect 3773 2597 3827 2603
rect 3773 2584 3779 2597
rect 3821 2584 3827 2597
rect 3725 2424 3731 2516
rect 3693 2417 3715 2423
rect 3533 2224 3539 2316
rect 3597 2304 3603 2336
rect 3613 2324 3619 2336
rect 3549 2143 3555 2276
rect 3533 2137 3555 2143
rect 3341 1843 3347 1956
rect 3373 1923 3379 2016
rect 3373 1917 3388 1923
rect 3421 1904 3427 2036
rect 3357 1864 3363 1896
rect 3325 1837 3347 1843
rect 3309 1623 3315 1696
rect 3325 1684 3331 1837
rect 3341 1784 3347 1796
rect 3389 1784 3395 1796
rect 3437 1784 3443 1996
rect 3469 1884 3475 2136
rect 3309 1617 3324 1623
rect 3325 1524 3331 1616
rect 3309 1504 3315 1516
rect 3357 1504 3363 1736
rect 3373 1724 3379 1736
rect 3421 1504 3427 1716
rect 3213 1484 3219 1496
rect 3149 1424 3155 1436
rect 3101 1144 3107 1336
rect 2637 1097 2652 1103
rect 2605 1064 2611 1096
rect 2573 744 2579 836
rect 2557 544 2563 656
rect 2589 583 2595 916
rect 2605 904 2611 1056
rect 2621 984 2627 1036
rect 2637 1004 2643 1097
rect 3117 1102 3123 1416
rect 3197 1404 3203 1476
rect 3229 1364 3235 1496
rect 3229 1324 3235 1336
rect 3213 1317 3228 1323
rect 3213 1104 3219 1317
rect 3245 1264 3251 1496
rect 3357 1484 3363 1496
rect 3373 1484 3379 1496
rect 3437 1484 3443 1496
rect 3277 1324 3283 1436
rect 3309 1344 3315 1476
rect 3341 1444 3347 1476
rect 3389 1444 3395 1456
rect 3373 1324 3379 1396
rect 3389 1244 3395 1316
rect 3229 1104 3235 1156
rect 3213 1084 3219 1096
rect 2909 1064 2915 1076
rect 3181 1064 3187 1076
rect 3245 1063 3251 1236
rect 3277 1104 3283 1236
rect 3229 1057 3251 1063
rect 2653 1037 2668 1043
rect 2621 844 2627 856
rect 2653 844 2659 1037
rect 2797 944 2803 1056
rect 2893 1037 2924 1043
rect 2893 1023 2899 1037
rect 2884 1017 2899 1023
rect 2813 926 2819 976
rect 2676 917 2691 923
rect 2877 924 2883 1016
rect 2938 1014 2950 1016
rect 2923 1006 2925 1014
rect 2933 1006 2935 1014
rect 2943 1006 2945 1014
rect 2953 1006 2955 1014
rect 2963 1006 2965 1014
rect 2938 1004 2950 1006
rect 2685 884 2691 917
rect 2621 724 2627 836
rect 2685 784 2691 836
rect 2893 824 2899 996
rect 2989 984 2995 1016
rect 3117 944 3123 1056
rect 3197 984 3203 1036
rect 3229 984 3235 1057
rect 3165 926 3171 976
rect 3197 924 3203 936
rect 2749 784 2755 816
rect 2621 684 2627 716
rect 2669 704 2675 716
rect 2573 577 2595 583
rect 2429 504 2435 536
rect 2420 297 2435 303
rect 2429 284 2435 297
rect 2317 203 2323 236
rect 2301 197 2323 203
rect 2285 124 2291 136
rect 2244 117 2259 123
rect 1933 104 1939 116
rect 2301 104 2307 197
rect 2349 184 2355 196
rect 2413 164 2419 236
rect 2429 224 2435 276
rect 2445 264 2451 536
rect 2461 304 2467 396
rect 2493 384 2499 476
rect 2509 384 2515 516
rect 2541 504 2547 516
rect 2573 404 2579 577
rect 2621 564 2627 676
rect 2653 544 2659 596
rect 2685 524 2691 776
rect 2717 524 2723 716
rect 2733 644 2739 776
rect 2781 724 2787 756
rect 2733 524 2739 636
rect 2749 624 2755 696
rect 2749 584 2755 616
rect 2781 544 2787 556
rect 2797 544 2803 656
rect 2829 543 2835 656
rect 2845 564 2851 676
rect 2861 664 2867 716
rect 2877 704 2883 736
rect 2893 684 2899 736
rect 2893 584 2899 656
rect 2909 644 2915 836
rect 3021 784 3027 916
rect 2941 664 2947 716
rect 3005 664 3011 716
rect 3101 704 3107 876
rect 3053 664 3059 696
rect 3085 664 3091 676
rect 3133 663 3139 836
rect 3197 784 3203 816
rect 3261 704 3267 876
rect 3325 702 3331 1036
rect 3357 964 3363 1076
rect 3405 984 3411 1436
rect 3421 1384 3427 1436
rect 3453 1324 3459 1776
rect 3469 1744 3475 1836
rect 3485 1724 3491 1876
rect 3501 1804 3507 1916
rect 3501 1764 3507 1776
rect 3517 1744 3523 2116
rect 3533 2104 3539 2137
rect 3549 2044 3555 2116
rect 3565 1964 3571 2156
rect 3597 2144 3603 2236
rect 3613 2184 3619 2316
rect 3693 2303 3699 2396
rect 3709 2383 3715 2417
rect 3709 2377 3731 2383
rect 3709 2324 3715 2356
rect 3693 2297 3715 2303
rect 3629 2284 3635 2296
rect 3661 2264 3667 2276
rect 3629 2184 3635 2236
rect 3661 2224 3667 2256
rect 3677 2184 3683 2296
rect 3709 2284 3715 2297
rect 3693 2164 3699 2276
rect 3725 2184 3731 2377
rect 3741 2344 3747 2556
rect 3757 2524 3763 2556
rect 3773 2444 3779 2476
rect 3773 2324 3779 2416
rect 3789 2343 3795 2576
rect 3837 2564 3843 2617
rect 3869 2584 3875 2756
rect 3901 2744 3907 2896
rect 3917 2884 3923 2897
rect 3901 2644 3907 2716
rect 3917 2604 3923 2696
rect 3949 2623 3955 2856
rect 3981 2784 3987 2936
rect 3965 2704 3971 2756
rect 3997 2684 4003 2936
rect 4029 2904 4035 3016
rect 4141 2984 4147 3076
rect 4301 3064 4307 3116
rect 4365 3104 4371 3176
rect 4324 3097 4339 3103
rect 4157 2964 4163 2976
rect 4084 2937 4099 2943
rect 4093 2923 4099 2937
rect 4125 2924 4131 2936
rect 4173 2924 4179 2996
rect 4093 2917 4108 2923
rect 4157 2903 4163 2916
rect 4157 2897 4188 2903
rect 4093 2744 4099 2896
rect 4109 2784 4115 2876
rect 4004 2677 4012 2683
rect 3981 2657 3996 2663
rect 3949 2617 3971 2623
rect 3805 2524 3811 2556
rect 3869 2544 3875 2556
rect 3885 2504 3891 2596
rect 3949 2584 3955 2596
rect 3901 2463 3907 2516
rect 3869 2457 3907 2463
rect 3869 2444 3875 2457
rect 3789 2337 3811 2343
rect 3757 2284 3763 2296
rect 3581 1904 3587 2016
rect 3549 1884 3555 1896
rect 3469 1684 3475 1716
rect 3469 1384 3475 1676
rect 3501 1504 3507 1676
rect 3549 1543 3555 1736
rect 3597 1724 3603 2136
rect 3613 1884 3619 1896
rect 3629 1844 3635 2096
rect 3725 2044 3731 2096
rect 3757 2044 3763 2276
rect 3773 2244 3779 2296
rect 3789 2184 3795 2316
rect 3805 2304 3811 2337
rect 3821 2304 3827 2396
rect 3901 2344 3907 2416
rect 3837 2184 3843 2276
rect 3853 2264 3859 2316
rect 3869 2244 3875 2316
rect 3885 2184 3891 2276
rect 3773 2144 3779 2176
rect 3837 2144 3843 2176
rect 3677 1984 3683 2036
rect 3533 1537 3555 1543
rect 3533 1524 3539 1537
rect 3549 1484 3555 1516
rect 3501 1444 3507 1476
rect 3517 1324 3523 1356
rect 3533 1344 3539 1476
rect 3565 1344 3571 1516
rect 3613 1504 3619 1676
rect 3597 1444 3603 1476
rect 3581 1344 3587 1436
rect 3565 1323 3571 1336
rect 3597 1324 3603 1416
rect 3613 1324 3619 1496
rect 3629 1424 3635 1816
rect 3645 1784 3651 1856
rect 3661 1844 3667 1916
rect 3693 1884 3699 1896
rect 3709 1884 3715 2036
rect 3677 1844 3683 1876
rect 3709 1784 3715 1856
rect 3725 1764 3731 1836
rect 3645 1684 3651 1718
rect 3677 1684 3683 1756
rect 3741 1724 3747 1876
rect 3757 1744 3763 1996
rect 3773 1884 3779 2116
rect 3789 2004 3795 2096
rect 3805 1884 3811 2036
rect 3869 1904 3875 1916
rect 3773 1784 3779 1856
rect 3805 1724 3811 1876
rect 3821 1844 3827 1896
rect 3869 1884 3875 1896
rect 3837 1864 3843 1876
rect 3837 1744 3843 1796
rect 3901 1784 3907 2336
rect 3917 2304 3923 2556
rect 3933 2544 3939 2556
rect 3965 2524 3971 2617
rect 3981 2584 3987 2657
rect 4029 2643 4035 2696
rect 4013 2637 4035 2643
rect 3981 2544 3987 2556
rect 3956 2497 3980 2503
rect 3997 2384 4003 2636
rect 4013 2564 4019 2637
rect 4061 2564 4067 2736
rect 4109 2703 4115 2736
rect 4157 2724 4163 2736
rect 4205 2724 4211 3036
rect 4100 2697 4115 2703
rect 4077 2604 4083 2676
rect 4157 2664 4163 2696
rect 4093 2584 4099 2596
rect 4013 2484 4019 2556
rect 4045 2524 4051 2556
rect 4077 2523 4083 2576
rect 4109 2564 4115 2656
rect 4125 2604 4131 2656
rect 4093 2544 4099 2556
rect 4077 2517 4115 2523
rect 3933 2304 3939 2316
rect 3965 2284 3971 2336
rect 3981 2304 3987 2336
rect 3997 2324 4003 2336
rect 3997 2264 4003 2296
rect 3933 2184 3939 2196
rect 3917 1904 3923 2116
rect 3917 1764 3923 1896
rect 3933 1864 3939 1916
rect 3949 1904 3955 2216
rect 3981 2144 3987 2176
rect 3965 2004 3971 2116
rect 3997 1963 4003 2176
rect 4013 2104 4019 2316
rect 4029 2224 4035 2516
rect 4045 2424 4051 2516
rect 4109 2504 4115 2517
rect 4093 2384 4099 2416
rect 4125 2383 4131 2576
rect 4141 2544 4147 2656
rect 4157 2503 4163 2516
rect 4157 2497 4188 2503
rect 4205 2424 4211 2656
rect 4221 2604 4227 2936
rect 4237 2924 4243 3036
rect 4301 2984 4307 2996
rect 4269 2924 4275 2956
rect 4333 2924 4339 3097
rect 4388 3077 4403 3083
rect 4365 3044 4371 3076
rect 4365 2983 4371 3036
rect 4397 2984 4403 3077
rect 4413 3064 4419 3176
rect 4413 3024 4419 3056
rect 4509 3043 4515 3296
rect 4541 3184 4547 3316
rect 4493 3037 4515 3043
rect 4413 2984 4419 3016
rect 4365 2977 4387 2983
rect 4365 2924 4371 2956
rect 4237 2744 4243 2916
rect 4317 2904 4323 2916
rect 4381 2904 4387 2977
rect 4221 2504 4227 2536
rect 4237 2524 4243 2736
rect 4253 2704 4259 2856
rect 4269 2704 4275 2856
rect 4333 2744 4339 2816
rect 4349 2784 4355 2876
rect 4413 2864 4419 2936
rect 4442 2814 4454 2816
rect 4427 2806 4429 2814
rect 4437 2806 4439 2814
rect 4447 2806 4449 2814
rect 4457 2806 4459 2814
rect 4467 2806 4469 2814
rect 4442 2804 4454 2806
rect 4381 2784 4387 2796
rect 4493 2784 4499 3037
rect 4541 2984 4547 3016
rect 4573 2984 4579 3276
rect 4605 3084 4611 3336
rect 4637 3326 4643 3336
rect 4605 3024 4611 3076
rect 4605 2984 4611 2996
rect 4509 2944 4515 2956
rect 4525 2944 4531 2956
rect 4541 2784 4547 2956
rect 4589 2804 4595 2956
rect 4605 2884 4611 2896
rect 4621 2784 4627 3236
rect 4685 3184 4691 3416
rect 4701 3344 4707 3476
rect 4733 3444 4739 3476
rect 4829 3404 4835 3476
rect 4861 3384 4867 3496
rect 4733 3084 4739 3196
rect 4781 3104 4787 3196
rect 4845 3184 4851 3296
rect 4877 3244 4883 3636
rect 4893 3584 4899 3757
rect 4909 3404 4915 3736
rect 4973 3704 4979 3776
rect 5021 3744 5027 3776
rect 5037 3744 5043 3856
rect 5053 3764 5059 3896
rect 5101 3884 5107 3896
rect 5085 3824 5091 3856
rect 5117 3804 5123 3896
rect 5069 3744 5075 3796
rect 4989 3584 4995 3656
rect 4925 3484 4931 3496
rect 4893 3084 4899 3316
rect 4708 3057 4723 3063
rect 4637 2904 4643 2956
rect 4669 2784 4675 2816
rect 4253 2664 4259 2696
rect 4285 2683 4291 2696
rect 4269 2677 4291 2683
rect 4253 2503 4259 2596
rect 4237 2497 4259 2503
rect 4109 2377 4131 2383
rect 4045 2264 4051 2296
rect 4077 2264 4083 2336
rect 4109 2284 4115 2377
rect 4125 2344 4131 2356
rect 4173 2284 4179 2296
rect 4157 2264 4163 2276
rect 4077 2184 4083 2236
rect 4109 2204 4115 2256
rect 4189 2244 4195 2376
rect 4109 2184 4115 2196
rect 4125 2164 4131 2236
rect 4093 2144 4099 2156
rect 4157 2144 4163 2216
rect 4221 2184 4227 2416
rect 4237 2404 4243 2497
rect 4253 2404 4259 2436
rect 4253 2263 4259 2356
rect 4269 2344 4275 2677
rect 4301 2664 4307 2676
rect 4285 2584 4291 2616
rect 4349 2503 4355 2696
rect 4413 2544 4419 2776
rect 4685 2764 4691 2936
rect 4717 2843 4723 3057
rect 4749 2964 4755 3016
rect 4765 2924 4771 3076
rect 4813 2984 4819 3056
rect 4717 2837 4739 2843
rect 4333 2497 4355 2503
rect 4269 2304 4275 2316
rect 4253 2257 4268 2263
rect 4189 2140 4195 2156
rect 4237 2144 4243 2216
rect 4253 2164 4259 2236
rect 4061 2084 4067 2096
rect 4029 2064 4035 2076
rect 3997 1957 4019 1963
rect 3972 1917 3996 1923
rect 4013 1904 4019 1957
rect 4029 1904 4035 2036
rect 4061 1984 4067 1996
rect 4077 1904 4083 1916
rect 3997 1864 4003 1896
rect 3981 1784 3987 1856
rect 4013 1784 4019 1816
rect 4045 1784 4051 1856
rect 4093 1784 4099 1916
rect 4029 1764 4035 1776
rect 4109 1763 4115 1916
rect 4125 1904 4131 1996
rect 4173 1944 4179 1956
rect 4205 1924 4211 2096
rect 4237 2024 4243 2116
rect 4221 1984 4227 2016
rect 4253 1984 4259 1996
rect 4212 1917 4220 1923
rect 4189 1864 4195 1896
rect 4093 1757 4115 1763
rect 3645 1584 3651 1616
rect 3565 1317 3587 1323
rect 3437 1244 3443 1296
rect 3565 1284 3571 1296
rect 3437 1124 3443 1236
rect 3485 1124 3491 1236
rect 3357 926 3363 936
rect 3389 924 3395 936
rect 3437 903 3443 1116
rect 3469 1084 3475 1096
rect 3501 1084 3507 1196
rect 3549 1104 3555 1196
rect 3565 1184 3571 1256
rect 3533 1084 3539 1096
rect 3453 1064 3459 1076
rect 3501 984 3507 996
rect 3485 964 3491 976
rect 3469 944 3475 956
rect 3453 924 3459 936
rect 3428 897 3443 903
rect 3437 724 3443 897
rect 3485 704 3491 936
rect 3549 924 3555 1076
rect 3533 884 3539 916
rect 3565 844 3571 1036
rect 3581 1024 3587 1317
rect 3645 1303 3651 1476
rect 3661 1444 3667 1516
rect 3693 1484 3699 1676
rect 3709 1624 3715 1696
rect 3709 1484 3715 1516
rect 3709 1424 3715 1436
rect 3677 1324 3683 1416
rect 3725 1363 3731 1636
rect 3773 1624 3779 1696
rect 3789 1503 3795 1656
rect 3821 1563 3827 1736
rect 3885 1624 3891 1696
rect 3901 1624 3907 1736
rect 3933 1724 3939 1736
rect 3812 1557 3827 1563
rect 3805 1524 3811 1556
rect 3837 1544 3843 1596
rect 3853 1543 3859 1556
rect 3853 1537 3891 1543
rect 3885 1524 3891 1537
rect 3789 1497 3811 1503
rect 3757 1444 3763 1476
rect 3773 1423 3779 1496
rect 3757 1417 3779 1423
rect 3716 1357 3731 1363
rect 3725 1324 3731 1357
rect 3636 1297 3651 1303
rect 3597 944 3603 1016
rect 3645 1004 3651 1236
rect 3661 983 3667 1296
rect 3741 1264 3747 1356
rect 3693 1124 3699 1236
rect 3757 1104 3763 1417
rect 3773 1384 3779 1396
rect 3789 1284 3795 1356
rect 3773 1103 3779 1236
rect 3773 1097 3788 1103
rect 3645 977 3667 983
rect 3613 924 3619 936
rect 3645 904 3651 977
rect 3677 924 3683 1076
rect 3805 1064 3811 1497
rect 3821 1384 3827 1476
rect 3853 1444 3859 1496
rect 3901 1463 3907 1576
rect 3917 1504 3923 1716
rect 3949 1604 3955 1716
rect 3965 1584 3971 1736
rect 3997 1644 4003 1696
rect 4013 1584 4019 1756
rect 4061 1683 4067 1756
rect 4045 1677 4067 1683
rect 3933 1504 3939 1576
rect 3917 1464 3923 1476
rect 3885 1457 3907 1463
rect 3869 1344 3875 1456
rect 3885 1340 3891 1457
rect 3901 1424 3907 1436
rect 3949 1384 3955 1576
rect 4045 1544 4051 1677
rect 3837 1264 3843 1316
rect 3869 1304 3875 1336
rect 3725 964 3731 996
rect 3757 944 3763 1036
rect 3773 924 3779 1016
rect 3805 984 3811 1056
rect 3837 983 3843 1216
rect 3853 1184 3859 1276
rect 3885 1143 3891 1332
rect 3949 1324 3955 1336
rect 3869 1137 3891 1143
rect 3869 1064 3875 1137
rect 3869 1044 3875 1056
rect 3853 1003 3859 1036
rect 3869 1024 3875 1036
rect 3853 997 3875 1003
rect 3837 977 3859 983
rect 3501 704 3507 756
rect 3133 657 3155 663
rect 2938 614 2950 616
rect 2923 606 2925 614
rect 2933 606 2935 614
rect 2943 606 2945 614
rect 2953 606 2955 614
rect 2963 606 2965 614
rect 2938 604 2950 606
rect 2845 544 2851 556
rect 2820 537 2835 543
rect 2797 524 2803 536
rect 2877 524 2883 556
rect 2861 517 2876 523
rect 2637 504 2643 516
rect 2749 504 2755 516
rect 2813 504 2819 516
rect 2605 344 2611 436
rect 2637 424 2643 496
rect 2477 283 2483 316
rect 2509 304 2515 336
rect 2637 304 2643 336
rect 2461 277 2483 283
rect 2461 184 2467 277
rect 2477 144 2483 256
rect 2493 184 2499 296
rect 2589 244 2595 276
rect 2669 264 2675 376
rect 2317 104 2323 136
rect 2525 124 2531 236
rect 2589 144 2595 196
rect 2685 164 2691 276
rect 2701 264 2707 436
rect 2717 304 2723 336
rect 2733 304 2739 316
rect 2765 284 2771 296
rect 2765 244 2771 276
rect 2813 184 2819 356
rect 2845 184 2851 256
rect 2861 204 2867 517
rect 2909 324 2915 476
rect 2877 224 2883 316
rect 2909 304 2915 316
rect 2925 304 2931 576
rect 3053 544 3059 636
rect 3133 544 3139 636
rect 3037 537 3052 543
rect 3012 317 3027 323
rect 2957 284 2963 296
rect 2938 214 2950 216
rect 2923 206 2925 214
rect 2933 206 2935 214
rect 2943 206 2945 214
rect 2953 206 2955 214
rect 2963 206 2965 214
rect 2938 204 2950 206
rect 2717 164 2723 176
rect 2765 164 2771 176
rect 2605 124 2611 156
rect 2637 124 2643 136
rect 2653 124 2659 136
rect 2813 124 2819 176
rect 2861 144 2867 196
rect 2989 163 2995 276
rect 3021 184 3027 317
rect 3037 203 3043 537
rect 3053 304 3059 396
rect 3117 364 3123 436
rect 3133 384 3139 536
rect 3149 524 3155 657
rect 3181 583 3187 696
rect 3172 577 3187 583
rect 3165 504 3171 576
rect 3101 324 3107 336
rect 3069 264 3075 276
rect 3037 197 3059 203
rect 3037 164 3043 176
rect 3053 164 3059 197
rect 3117 184 3123 256
rect 2980 157 2995 163
rect 2909 124 2915 136
rect 3053 124 3059 156
rect 3133 124 3139 316
rect 3149 264 3155 276
rect 3165 264 3171 376
rect 3229 304 3235 656
rect 3261 544 3267 696
rect 3485 684 3491 696
rect 3421 524 3427 536
rect 3469 524 3475 636
rect 3485 526 3491 596
rect 3581 544 3587 836
rect 3645 824 3651 896
rect 3597 523 3603 816
rect 3661 783 3667 836
rect 3645 777 3667 783
rect 3645 702 3651 777
rect 3677 684 3683 916
rect 3709 684 3715 856
rect 3725 844 3731 916
rect 3757 724 3763 816
rect 3588 517 3603 523
rect 3357 404 3363 436
rect 3549 384 3555 436
rect 3149 124 3155 236
rect 3197 144 3203 236
rect 3229 124 3235 256
rect 3245 184 3251 196
rect 3341 164 3347 276
rect 3373 264 3379 356
rect 3405 284 3411 336
rect 3373 126 3379 176
rect 3485 164 3491 276
rect 3501 124 3507 376
rect 3661 304 3667 316
rect 3677 124 3683 496
rect 3709 304 3715 536
rect 3773 404 3779 916
rect 3789 884 3795 936
rect 3821 924 3827 936
rect 3837 904 3843 936
rect 3805 724 3811 836
rect 3853 784 3859 977
rect 3869 923 3875 997
rect 3885 964 3891 1116
rect 3917 1084 3923 1296
rect 3933 1224 3939 1296
rect 3965 1284 3971 1356
rect 3981 1304 3987 1436
rect 3997 1364 4003 1536
rect 4093 1523 4099 1757
rect 4205 1763 4211 1876
rect 4221 1784 4227 1916
rect 4269 1884 4275 2256
rect 4285 2203 4291 2436
rect 4301 2244 4307 2256
rect 4285 2197 4307 2203
rect 4301 2184 4307 2197
rect 4317 2084 4323 2236
rect 4333 2224 4339 2497
rect 4413 2464 4419 2536
rect 4461 2504 4467 2656
rect 4442 2414 4454 2416
rect 4427 2406 4429 2414
rect 4437 2406 4439 2414
rect 4447 2406 4449 2414
rect 4457 2406 4459 2414
rect 4467 2406 4469 2414
rect 4442 2404 4454 2406
rect 4397 2344 4403 2396
rect 4493 2364 4499 2736
rect 4653 2724 4659 2756
rect 4733 2724 4739 2837
rect 4509 2584 4515 2676
rect 4525 2544 4531 2656
rect 4541 2584 4547 2656
rect 4397 2284 4403 2296
rect 4365 2183 4371 2256
rect 4365 2177 4387 2183
rect 4365 2144 4371 2156
rect 4349 2124 4355 2136
rect 4333 1984 4339 2116
rect 4333 1964 4339 1976
rect 4285 1924 4291 1956
rect 4324 1877 4339 1883
rect 4237 1784 4243 1856
rect 4253 1764 4259 1856
rect 4269 1843 4275 1856
rect 4269 1837 4291 1843
rect 4285 1764 4291 1837
rect 4333 1784 4339 1877
rect 4205 1757 4227 1763
rect 4125 1744 4131 1756
rect 4109 1564 4115 1696
rect 4125 1584 4131 1716
rect 4157 1524 4163 1656
rect 4093 1517 4115 1523
rect 4013 1384 4019 1496
rect 4029 1444 4035 1516
rect 4077 1464 4083 1476
rect 4093 1444 4099 1476
rect 4013 1364 4019 1376
rect 4013 1344 4019 1356
rect 3981 1184 3987 1236
rect 4029 1163 4035 1356
rect 4045 1344 4051 1376
rect 4109 1364 4115 1517
rect 4141 1483 4147 1516
rect 4125 1477 4147 1483
rect 4077 1324 4083 1356
rect 4077 1304 4083 1316
rect 4013 1157 4035 1163
rect 3949 1084 3955 1136
rect 3981 1104 3987 1136
rect 3901 944 3907 1036
rect 3917 1004 3923 1076
rect 3933 984 3939 1076
rect 3965 1063 3971 1096
rect 3997 1064 4003 1136
rect 4013 1084 4019 1157
rect 3949 1057 3971 1063
rect 3949 984 3955 1057
rect 3933 964 3939 976
rect 3869 917 3884 923
rect 3917 923 3923 956
rect 3965 944 3971 956
rect 3908 917 3923 923
rect 3869 824 3875 856
rect 3869 724 3875 816
rect 3949 724 3955 836
rect 3805 684 3811 696
rect 3789 604 3795 636
rect 3821 624 3827 696
rect 3869 663 3875 716
rect 3933 704 3939 716
rect 3965 704 3971 896
rect 3981 824 3987 1056
rect 3997 944 4003 1056
rect 4045 1044 4051 1096
rect 4013 904 4019 916
rect 3901 664 3907 696
rect 3917 684 3923 696
rect 3997 664 4003 696
rect 4029 664 4035 996
rect 4045 984 4051 1036
rect 4061 784 4067 1056
rect 4077 743 4083 1276
rect 4093 1184 4099 1296
rect 4109 1284 4115 1356
rect 4109 1184 4115 1256
rect 4125 1163 4131 1477
rect 4157 1384 4163 1516
rect 4173 1364 4179 1736
rect 4205 1664 4211 1736
rect 4189 1657 4204 1663
rect 4189 1484 4195 1657
rect 4189 1464 4195 1476
rect 4109 1157 4131 1163
rect 4109 1124 4115 1157
rect 4109 1004 4115 1096
rect 4125 984 4131 1116
rect 4141 1084 4147 1316
rect 4157 1204 4163 1316
rect 4173 1244 4179 1356
rect 4189 1344 4195 1416
rect 4205 1263 4211 1476
rect 4221 1443 4227 1757
rect 4349 1763 4355 2096
rect 4365 1923 4371 2096
rect 4381 2024 4387 2177
rect 4413 2084 4419 2296
rect 4461 2184 4467 2276
rect 4493 2184 4499 2336
rect 4509 2164 4515 2496
rect 4525 2484 4531 2536
rect 4541 2463 4547 2556
rect 4557 2483 4563 2656
rect 4573 2604 4579 2636
rect 4589 2564 4595 2676
rect 4557 2477 4572 2483
rect 4541 2457 4563 2463
rect 4525 2384 4531 2456
rect 4541 2404 4547 2436
rect 4557 2364 4563 2457
rect 4589 2384 4595 2556
rect 4605 2504 4611 2716
rect 4621 2483 4627 2496
rect 4637 2484 4643 2616
rect 4685 2584 4691 2676
rect 4701 2564 4707 2676
rect 4717 2624 4723 2636
rect 4733 2584 4739 2716
rect 4749 2684 4755 2856
rect 4845 2704 4851 2776
rect 4717 2563 4723 2576
rect 4717 2557 4739 2563
rect 4733 2544 4739 2557
rect 4653 2504 4659 2536
rect 4612 2477 4627 2483
rect 4669 2384 4675 2416
rect 4541 2183 4547 2356
rect 4621 2344 4627 2356
rect 4557 2284 4563 2296
rect 4637 2284 4643 2296
rect 4685 2244 4691 2516
rect 4701 2384 4707 2536
rect 4717 2404 4723 2536
rect 4724 2337 4739 2343
rect 4733 2264 4739 2337
rect 4749 2324 4755 2676
rect 4781 2584 4787 2676
rect 4813 2544 4819 2556
rect 4829 2544 4835 2616
rect 4541 2177 4556 2183
rect 4477 2104 4483 2156
rect 4541 2144 4547 2156
rect 4388 2017 4403 2023
rect 4397 1984 4403 2017
rect 4442 2014 4454 2016
rect 4427 2006 4429 2014
rect 4437 2006 4439 2014
rect 4447 2006 4449 2014
rect 4457 2006 4459 2014
rect 4467 2006 4469 2014
rect 4442 2004 4454 2006
rect 4381 1943 4387 1976
rect 4381 1937 4396 1943
rect 4365 1917 4380 1923
rect 4397 1897 4412 1903
rect 4365 1784 4371 1816
rect 4333 1757 4355 1763
rect 4237 1484 4243 1756
rect 4221 1437 4243 1443
rect 4189 1257 4211 1263
rect 4141 1064 4147 1076
rect 4093 964 4099 976
rect 4125 964 4131 976
rect 4093 904 4099 916
rect 4125 904 4131 916
rect 4141 883 4147 896
rect 4132 877 4147 883
rect 4157 784 4163 1156
rect 4173 1084 4179 1116
rect 4189 1084 4195 1257
rect 4205 1104 4211 1236
rect 4221 1184 4227 1276
rect 4237 1184 4243 1437
rect 4253 1424 4259 1756
rect 4317 1744 4323 1756
rect 4333 1723 4339 1757
rect 4317 1717 4339 1723
rect 4317 1584 4323 1717
rect 4397 1703 4403 1897
rect 4349 1697 4403 1703
rect 4349 1644 4355 1697
rect 4445 1644 4451 1976
rect 4461 1764 4467 1976
rect 4493 1884 4499 2116
rect 4509 1984 4515 2036
rect 4573 1984 4579 2236
rect 4749 2224 4755 2276
rect 4605 2104 4611 2136
rect 4621 2104 4627 2196
rect 4765 2184 4771 2516
rect 4781 2444 4787 2476
rect 4813 2304 4819 2316
rect 4797 2264 4803 2296
rect 4829 2204 4835 2236
rect 4644 2157 4739 2163
rect 4733 2144 4739 2157
rect 4845 2144 4851 2696
rect 4861 2584 4867 3076
rect 4893 2944 4899 3076
rect 4925 3023 4931 3436
rect 4957 3364 4963 3376
rect 4973 3344 4979 3396
rect 5005 3384 5011 3496
rect 5021 3464 5027 3496
rect 5037 3384 5043 3496
rect 5053 3484 5059 3716
rect 5085 3664 5091 3796
rect 5149 3764 5155 4196
rect 5197 4184 5203 4237
rect 5229 4164 5235 4476
rect 5261 4344 5267 4556
rect 5293 4504 5299 4557
rect 5261 4304 5267 4336
rect 5229 4124 5235 4136
rect 5245 4123 5251 4296
rect 5261 4277 5276 4283
rect 5261 4144 5267 4277
rect 5293 4244 5299 4296
rect 5309 4284 5315 4456
rect 5325 4304 5331 4416
rect 5341 4344 5347 4696
rect 5357 4604 5363 4636
rect 5373 4524 5379 4716
rect 5453 4704 5459 4916
rect 5485 4764 5491 4896
rect 5485 4604 5491 4694
rect 5517 4684 5523 4936
rect 5549 4744 5555 4956
rect 5565 4864 5571 5076
rect 5581 4864 5587 4916
rect 5597 4904 5603 5076
rect 5645 4964 5651 5056
rect 5597 4784 5603 4816
rect 5565 4704 5571 4756
rect 5389 4524 5395 4596
rect 5437 4524 5443 4576
rect 5469 4524 5475 4556
rect 5501 4524 5507 4616
rect 5533 4584 5539 4596
rect 5549 4544 5555 4616
rect 5581 4564 5587 4776
rect 5661 4764 5667 5216
rect 5725 5124 5731 5216
rect 5773 5123 5779 5136
rect 5773 5117 5795 5123
rect 5789 5104 5795 5117
rect 5677 4984 5683 5056
rect 5693 5004 5699 5096
rect 5709 5024 5715 5036
rect 5741 4944 5747 5036
rect 5757 4924 5763 4936
rect 5773 4924 5779 5096
rect 5805 5083 5811 5136
rect 5837 5104 5843 5116
rect 5853 5103 5859 5276
rect 5869 5124 5875 5236
rect 5853 5097 5875 5103
rect 5869 5084 5875 5097
rect 5796 5077 5811 5083
rect 5853 5044 5859 5076
rect 5789 4924 5795 5016
rect 5805 4944 5811 5036
rect 5901 5024 5907 5256
rect 5917 5104 5923 5316
rect 6125 5184 6131 5196
rect 6157 5164 6163 5336
rect 6269 5324 6275 5336
rect 6317 5324 6323 5356
rect 6365 5324 6371 5336
rect 6413 5324 6419 5356
rect 6493 5344 6499 5376
rect 6797 5344 6803 5376
rect 6461 5324 6467 5336
rect 6285 5224 6291 5316
rect 6381 5303 6387 5316
rect 6372 5297 6387 5303
rect 5933 5044 5939 5116
rect 5997 5104 6003 5156
rect 6013 5104 6019 5136
rect 6157 5104 6163 5136
rect 6109 5064 6115 5096
rect 6173 5044 6179 5096
rect 6221 5064 6227 5116
rect 6285 5104 6291 5216
rect 6333 5184 6339 5236
rect 6333 5144 6339 5156
rect 6301 5124 6307 5136
rect 6269 5084 6275 5096
rect 5946 5014 5958 5016
rect 5931 5006 5933 5014
rect 5941 5006 5943 5014
rect 5951 5006 5953 5014
rect 5961 5006 5963 5014
rect 5971 5006 5973 5014
rect 5946 5004 5958 5006
rect 5677 4743 5683 4836
rect 5668 4737 5683 4743
rect 5693 4704 5699 4856
rect 5629 4684 5635 4696
rect 5725 4684 5731 4916
rect 5741 4744 5747 4916
rect 5757 4844 5763 4856
rect 5757 4683 5763 4836
rect 5789 4784 5795 4836
rect 5805 4764 5811 4936
rect 5853 4924 5859 4996
rect 5885 4924 5891 4976
rect 6029 4924 6035 4936
rect 6077 4924 6083 4996
rect 6189 4944 6195 4976
rect 5773 4704 5779 4736
rect 5757 4677 5779 4683
rect 5581 4524 5587 4556
rect 5613 4524 5619 4676
rect 5725 4664 5731 4676
rect 5357 4504 5363 4516
rect 5565 4503 5571 4516
rect 5565 4497 5587 4503
rect 5405 4424 5411 4436
rect 5501 4384 5507 4456
rect 5565 4304 5571 4336
rect 5277 4124 5283 4156
rect 5293 4144 5299 4156
rect 5245 4117 5267 4123
rect 5229 4097 5244 4103
rect 5197 3904 5203 4036
rect 5229 3924 5235 4097
rect 5261 4044 5267 4117
rect 5213 3904 5219 3916
rect 5165 3804 5171 3876
rect 5181 3824 5187 3856
rect 5197 3764 5203 3896
rect 5229 3864 5235 3916
rect 5245 3844 5251 3976
rect 5277 3903 5283 4116
rect 5309 4104 5315 4276
rect 5341 4124 5347 4256
rect 5357 4204 5363 4296
rect 5421 4264 5427 4296
rect 5389 4204 5395 4256
rect 5469 4224 5475 4296
rect 5533 4284 5539 4296
rect 5549 4244 5555 4276
rect 5581 4243 5587 4497
rect 5613 4344 5619 4436
rect 5597 4264 5603 4296
rect 5613 4244 5619 4276
rect 5581 4237 5603 4243
rect 5357 4184 5363 4196
rect 5389 4104 5395 4116
rect 5309 4084 5315 4096
rect 5293 3944 5299 4076
rect 5268 3897 5283 3903
rect 5101 3724 5107 3736
rect 5117 3704 5123 3756
rect 5149 3724 5155 3756
rect 5213 3744 5219 3836
rect 5261 3824 5267 3896
rect 5277 3864 5283 3876
rect 5101 3484 5107 3496
rect 5133 3484 5139 3536
rect 5085 3364 5091 3376
rect 5149 3364 5155 3716
rect 5165 3704 5171 3736
rect 5229 3724 5235 3816
rect 5277 3784 5283 3816
rect 5229 3504 5235 3716
rect 5277 3704 5283 3756
rect 5293 3664 5299 3756
rect 5325 3744 5331 3916
rect 5421 3884 5427 3894
rect 5485 3884 5491 3936
rect 5501 3904 5507 4236
rect 5517 4064 5523 4116
rect 5533 3984 5539 4196
rect 5565 4144 5571 4176
rect 5597 4144 5603 4237
rect 5613 4164 5619 4196
rect 5597 3924 5603 4136
rect 5453 3864 5459 3876
rect 5341 3744 5347 3816
rect 5421 3784 5427 3796
rect 5485 3784 5491 3836
rect 5325 3724 5331 3736
rect 5373 3717 5388 3723
rect 5341 3703 5347 3716
rect 5325 3697 5347 3703
rect 5325 3684 5331 3697
rect 5373 3584 5379 3717
rect 5405 3704 5411 3736
rect 5501 3724 5507 3836
rect 5517 3824 5523 3916
rect 5533 3784 5539 3876
rect 5565 3724 5571 3816
rect 5421 3504 5427 3556
rect 5069 3344 5075 3356
rect 4989 3264 4995 3316
rect 5037 3264 5043 3296
rect 5117 3284 5123 3316
rect 5165 3284 5171 3336
rect 5181 3324 5187 3396
rect 5213 3344 5219 3496
rect 5293 3424 5299 3496
rect 5341 3384 5347 3496
rect 5389 3484 5395 3496
rect 5405 3464 5411 3496
rect 5421 3404 5427 3496
rect 5437 3484 5443 3496
rect 5133 3124 5139 3256
rect 4909 3017 4931 3023
rect 4877 2544 4883 2596
rect 4893 2584 4899 2916
rect 4909 2784 4915 3017
rect 5021 2944 5027 2956
rect 5021 2864 5027 2936
rect 5101 2924 5107 2996
rect 5117 2903 5123 3076
rect 5165 3064 5171 3076
rect 5165 3044 5171 3056
rect 5197 2984 5203 3096
rect 5245 2944 5251 3276
rect 5437 3204 5443 3476
rect 5453 3464 5459 3716
rect 5517 3704 5523 3716
rect 5533 3704 5539 3716
rect 5581 3644 5587 3736
rect 5629 3684 5635 4636
rect 5661 4584 5667 4636
rect 5661 4524 5667 4576
rect 5693 4544 5699 4596
rect 5725 4584 5731 4616
rect 5773 4584 5779 4677
rect 5789 4664 5795 4756
rect 5821 4724 5827 4916
rect 5837 4904 5843 4916
rect 5821 4584 5827 4696
rect 5837 4563 5843 4696
rect 5853 4584 5859 4916
rect 6093 4864 6099 4936
rect 6045 4824 6051 4836
rect 6109 4824 6115 4916
rect 6157 4884 6163 4936
rect 5917 4784 5923 4796
rect 5901 4704 5907 4756
rect 6077 4723 6083 4736
rect 6077 4717 6099 4723
rect 5965 4704 5971 4716
rect 5997 4624 6003 4696
rect 5946 4614 5958 4616
rect 5931 4606 5933 4614
rect 5941 4606 5943 4614
rect 5951 4606 5953 4614
rect 5961 4606 5963 4614
rect 5971 4606 5973 4614
rect 5946 4604 5958 4606
rect 5837 4557 5859 4563
rect 5709 4524 5715 4536
rect 5757 4524 5763 4556
rect 5645 4324 5651 4516
rect 5805 4504 5811 4516
rect 5661 4243 5667 4456
rect 5805 4384 5811 4496
rect 5821 4424 5827 4516
rect 5837 4344 5843 4416
rect 5677 4324 5683 4336
rect 5709 4304 5715 4336
rect 5773 4304 5779 4316
rect 5709 4284 5715 4296
rect 5741 4284 5747 4296
rect 5725 4264 5731 4276
rect 5645 4237 5667 4243
rect 5645 3843 5651 4237
rect 5661 4104 5667 4156
rect 5725 4144 5731 4236
rect 5693 4104 5699 4116
rect 5661 4084 5667 4096
rect 5709 4084 5715 4136
rect 5725 4124 5731 4136
rect 5757 4123 5763 4196
rect 5757 4117 5772 4123
rect 5789 4084 5795 4276
rect 5821 4163 5827 4316
rect 5853 4244 5859 4557
rect 5869 4524 5875 4536
rect 5901 4504 5907 4596
rect 6013 4584 6019 4676
rect 6029 4564 6035 4656
rect 5981 4524 5987 4536
rect 5917 4284 5923 4436
rect 5981 4403 5987 4516
rect 6029 4464 6035 4556
rect 6045 4504 6051 4596
rect 6061 4564 6067 4716
rect 6093 4704 6099 4717
rect 6141 4704 6147 4796
rect 6173 4724 6179 4936
rect 6205 4924 6211 4956
rect 6269 4924 6275 5036
rect 6285 4944 6291 4996
rect 6349 4944 6355 4996
rect 6365 4944 6371 5296
rect 6477 5284 6483 5316
rect 6573 5304 6579 5316
rect 6413 5064 6419 5096
rect 6461 5084 6467 5116
rect 6525 5084 6531 5096
rect 6461 5024 6467 5076
rect 6493 5044 6499 5056
rect 6493 5023 6499 5036
rect 6477 5017 6499 5023
rect 6333 4924 6339 4936
rect 6429 4924 6435 4976
rect 6461 4944 6467 4956
rect 6445 4924 6451 4936
rect 6477 4924 6483 5017
rect 6525 4924 6531 4976
rect 6541 4924 6547 5276
rect 6573 5103 6579 5236
rect 6589 5224 6595 5336
rect 6717 5284 6723 5316
rect 6637 5124 6643 5136
rect 6765 5104 6771 5336
rect 6925 5326 6931 5396
rect 7053 5384 7059 5396
rect 7197 5377 7212 5383
rect 6989 5364 6995 5376
rect 7197 5364 7203 5377
rect 7197 5344 7203 5356
rect 6829 5104 6835 5136
rect 6573 5097 6588 5103
rect 6557 4964 6563 4996
rect 6589 4983 6595 5096
rect 6765 5084 6771 5096
rect 6909 5084 6915 5096
rect 6957 5084 6963 5336
rect 7165 5324 7171 5336
rect 6637 4984 6643 5076
rect 6797 5004 6803 5036
rect 6589 4977 6611 4983
rect 6605 4924 6611 4977
rect 6941 4964 6947 4976
rect 6989 4944 6995 4956
rect 6276 4917 6291 4923
rect 6285 4844 6291 4917
rect 6301 4864 6307 4896
rect 6077 4524 6083 4696
rect 6093 4664 6099 4676
rect 6061 4504 6067 4516
rect 5981 4397 6003 4403
rect 5869 4264 5875 4276
rect 5805 4157 5827 4163
rect 5805 4124 5811 4157
rect 5821 4103 5827 4136
rect 5837 4124 5843 4196
rect 5853 4144 5859 4216
rect 5885 4164 5891 4276
rect 5901 4163 5907 4276
rect 5946 4214 5958 4216
rect 5931 4206 5933 4214
rect 5941 4206 5943 4214
rect 5951 4206 5953 4214
rect 5961 4206 5963 4214
rect 5971 4206 5973 4214
rect 5946 4204 5958 4206
rect 5901 4157 5923 4163
rect 5876 4117 5884 4123
rect 5901 4103 5907 4136
rect 5821 4097 5907 4103
rect 5789 4044 5795 4076
rect 5917 3984 5923 4157
rect 5933 4124 5939 4156
rect 5661 3902 5667 3936
rect 5725 3884 5731 3976
rect 5693 3864 5699 3876
rect 5757 3864 5763 3916
rect 5773 3884 5779 3936
rect 5693 3844 5699 3856
rect 5645 3837 5667 3843
rect 5645 3744 5651 3776
rect 5645 3664 5651 3716
rect 5581 3584 5587 3636
rect 5533 3484 5539 3496
rect 5485 3464 5491 3476
rect 5453 3424 5459 3436
rect 5389 3104 5395 3136
rect 5453 3123 5459 3136
rect 5437 3117 5459 3123
rect 5437 3104 5443 3117
rect 5261 2984 5267 2996
rect 5293 2984 5299 3096
rect 5293 2964 5299 2976
rect 5229 2924 5235 2936
rect 5245 2924 5251 2936
rect 5229 2904 5235 2916
rect 5101 2897 5123 2903
rect 5101 2744 5107 2897
rect 5229 2864 5235 2896
rect 5309 2844 5315 2976
rect 5341 2904 5347 2916
rect 5069 2702 5075 2716
rect 4909 2677 4924 2683
rect 4909 2524 4915 2677
rect 4957 2644 4963 2676
rect 4925 2504 4931 2636
rect 4941 2624 4947 2636
rect 5005 2544 5011 2556
rect 4605 1964 4611 2096
rect 4525 1864 4531 1896
rect 4541 1864 4547 1956
rect 4541 1763 4547 1856
rect 4541 1757 4556 1763
rect 4525 1724 4531 1756
rect 4461 1644 4467 1716
rect 4525 1704 4531 1716
rect 4381 1584 4387 1636
rect 4269 1544 4275 1576
rect 4292 1497 4307 1503
rect 4269 1104 4275 1296
rect 4301 1184 4307 1497
rect 4285 1124 4291 1176
rect 4196 1057 4211 1063
rect 4189 944 4195 1036
rect 4077 737 4099 743
rect 3853 657 3875 663
rect 3837 644 3843 656
rect 3853 563 3859 657
rect 3869 564 3875 636
rect 3901 564 3907 596
rect 3981 584 3987 656
rect 4045 604 4051 716
rect 4077 564 4083 656
rect 3844 557 3859 563
rect 3917 504 3923 556
rect 3949 524 3955 536
rect 3933 504 3939 516
rect 3796 297 3811 303
rect 3709 144 3715 296
rect 3789 264 3795 276
rect 3805 264 3811 297
rect 3853 284 3859 396
rect 3869 324 3875 436
rect 3917 384 3923 496
rect 4013 484 4019 496
rect 3757 184 3763 256
rect 3837 244 3843 256
rect 3821 184 3827 236
rect 3853 204 3859 276
rect 3908 257 3923 263
rect 3725 144 3731 156
rect 3853 124 3859 176
rect 3917 164 3923 257
rect 3933 244 3939 256
rect 3933 204 3939 236
rect 3949 184 3955 356
rect 4045 324 4051 556
rect 4093 384 4099 737
rect 4125 724 4131 736
rect 4173 704 4179 936
rect 4189 764 4195 936
rect 4205 924 4211 1057
rect 4221 824 4227 1096
rect 4237 984 4243 996
rect 4285 984 4291 1076
rect 4253 964 4259 976
rect 4285 964 4291 976
rect 4317 944 4323 1236
rect 4333 1144 4339 1536
rect 4365 1524 4371 1576
rect 4397 1563 4403 1636
rect 4442 1614 4454 1616
rect 4427 1606 4429 1614
rect 4437 1606 4439 1614
rect 4447 1606 4449 1614
rect 4457 1606 4459 1614
rect 4467 1606 4469 1614
rect 4442 1604 4454 1606
rect 4493 1564 4499 1596
rect 4509 1564 4515 1696
rect 4381 1557 4403 1563
rect 4349 1304 4355 1496
rect 4365 1304 4371 1336
rect 4381 1243 4387 1557
rect 4429 1244 4435 1516
rect 4509 1464 4515 1476
rect 4509 1324 4515 1356
rect 4381 1237 4403 1243
rect 4349 1144 4355 1216
rect 4365 903 4371 1116
rect 4349 897 4371 903
rect 4237 784 4243 896
rect 4253 784 4259 816
rect 4269 764 4275 836
rect 4317 784 4323 896
rect 4349 784 4355 897
rect 4221 724 4227 736
rect 4237 704 4243 756
rect 4292 717 4307 723
rect 4109 664 4115 676
rect 4157 644 4163 696
rect 4109 384 4115 616
rect 4205 584 4211 616
rect 4221 584 4227 676
rect 4301 664 4307 717
rect 4365 684 4371 856
rect 4397 784 4403 1237
rect 4442 1214 4454 1216
rect 4427 1206 4429 1214
rect 4437 1206 4439 1214
rect 4447 1206 4449 1214
rect 4457 1206 4459 1214
rect 4467 1206 4469 1214
rect 4442 1204 4454 1206
rect 4429 1164 4435 1176
rect 4493 1144 4499 1216
rect 4509 1204 4515 1316
rect 4509 1104 4515 1196
rect 4525 1184 4531 1376
rect 4541 1264 4547 1636
rect 4557 1584 4563 1656
rect 4573 1484 4579 1636
rect 4589 1524 4595 1916
rect 4605 1864 4611 1876
rect 4621 1864 4627 1876
rect 4621 1744 4627 1756
rect 4589 1424 4595 1496
rect 4541 1184 4547 1236
rect 4557 1184 4563 1416
rect 4413 926 4419 976
rect 4445 944 4451 1096
rect 4573 1064 4579 1318
rect 4605 1284 4611 1716
rect 4621 1544 4627 1676
rect 4637 1584 4643 2116
rect 4653 1944 4659 2136
rect 4701 2044 4707 2116
rect 4669 1784 4675 1916
rect 4717 1864 4723 2116
rect 4781 1944 4787 2056
rect 4797 1984 4803 2096
rect 4861 1984 4867 2456
rect 4909 2424 4915 2496
rect 4957 2323 4963 2476
rect 4941 2317 4963 2323
rect 4941 2184 4947 2317
rect 4957 2224 4963 2294
rect 4877 2124 4883 2136
rect 4973 2084 4979 2136
rect 4733 1897 4748 1903
rect 4669 1744 4675 1776
rect 4685 1704 4691 1756
rect 4621 1484 4627 1516
rect 4621 1184 4627 1256
rect 4653 1144 4659 1536
rect 4685 1364 4691 1636
rect 4717 1584 4723 1676
rect 4733 1563 4739 1897
rect 4804 1897 4819 1903
rect 4749 1584 4755 1856
rect 4765 1664 4771 1696
rect 4813 1584 4819 1897
rect 4829 1764 4835 1956
rect 4845 1884 4851 1896
rect 4877 1863 4883 2036
rect 4909 1984 4915 2036
rect 4877 1857 4899 1863
rect 4845 1784 4851 1796
rect 4893 1764 4899 1857
rect 4925 1764 4931 2076
rect 4973 2024 4979 2076
rect 4989 2004 4995 2276
rect 5021 2264 5027 2616
rect 5101 2524 5107 2736
rect 5053 2344 5059 2476
rect 5101 2364 5107 2496
rect 5133 2464 5139 2676
rect 5165 2504 5171 2696
rect 5181 2584 5187 2716
rect 5229 2704 5235 2716
rect 5197 2684 5203 2696
rect 5197 2544 5203 2616
rect 5213 2544 5219 2656
rect 5229 2543 5235 2696
rect 5252 2637 5267 2643
rect 5229 2537 5251 2543
rect 5133 2357 5148 2363
rect 5053 2317 5084 2323
rect 5053 2304 5059 2317
rect 5085 2284 5091 2296
rect 5133 2284 5139 2357
rect 5149 2324 5155 2356
rect 5069 2244 5075 2276
rect 5117 2184 5123 2216
rect 5069 2124 5075 2136
rect 5005 2104 5011 2116
rect 5069 2044 5075 2116
rect 5101 2064 5107 2136
rect 5165 2124 5171 2496
rect 5197 2404 5203 2536
rect 5181 2284 5187 2296
rect 5197 2284 5203 2336
rect 5213 2284 5219 2296
rect 5181 2164 5187 2196
rect 5181 2124 5187 2156
rect 5245 2143 5251 2537
rect 5261 2383 5267 2637
rect 5277 2524 5283 2576
rect 5325 2524 5331 2776
rect 5341 2704 5347 2896
rect 5357 2884 5363 3096
rect 5389 2784 5395 3036
rect 5437 2944 5443 3036
rect 5453 3004 5459 3076
rect 5469 2944 5475 3336
rect 5533 3284 5539 3476
rect 5565 3424 5571 3456
rect 5581 3344 5587 3536
rect 5629 3444 5635 3496
rect 5597 3364 5603 3436
rect 5565 3337 5580 3343
rect 5565 3304 5571 3337
rect 5597 3264 5603 3316
rect 5645 3264 5651 3296
rect 5661 3284 5667 3837
rect 5757 3824 5763 3856
rect 5677 3724 5683 3736
rect 5677 3504 5683 3596
rect 5693 3564 5699 3736
rect 5709 3564 5715 3716
rect 5725 3703 5731 3716
rect 5725 3697 5740 3703
rect 5789 3544 5795 3976
rect 5805 3864 5811 3896
rect 5837 3884 5843 3896
rect 5837 3704 5843 3876
rect 5677 3363 5683 3496
rect 5693 3444 5699 3496
rect 5709 3484 5715 3496
rect 5709 3423 5715 3476
rect 5789 3464 5795 3496
rect 5805 3484 5811 3496
rect 5693 3417 5715 3423
rect 5693 3384 5699 3417
rect 5725 3384 5731 3436
rect 5677 3357 5699 3363
rect 5677 3284 5683 3336
rect 5645 3184 5651 3196
rect 5677 3184 5683 3256
rect 5693 3224 5699 3357
rect 5789 3326 5795 3356
rect 5725 3304 5731 3316
rect 5517 3104 5523 3116
rect 5613 3104 5619 3156
rect 5709 3104 5715 3256
rect 5725 3143 5731 3296
rect 5725 3137 5747 3143
rect 5565 3084 5571 3096
rect 5597 3077 5612 3083
rect 5485 3044 5491 3056
rect 5581 3044 5587 3056
rect 5437 2764 5443 2916
rect 5437 2704 5443 2756
rect 5373 2664 5379 2694
rect 5469 2684 5475 2936
rect 5501 2926 5507 2936
rect 5485 2704 5491 2736
rect 5485 2664 5491 2696
rect 5501 2684 5507 2696
rect 5373 2524 5379 2616
rect 5437 2584 5443 2656
rect 5469 2643 5475 2656
rect 5469 2637 5491 2643
rect 5453 2564 5459 2636
rect 5261 2377 5276 2383
rect 5277 2304 5283 2376
rect 5309 2324 5315 2516
rect 5389 2484 5395 2516
rect 5405 2504 5411 2516
rect 5405 2464 5411 2496
rect 5421 2464 5427 2536
rect 5293 2284 5299 2296
rect 5229 2137 5251 2143
rect 5229 2124 5235 2137
rect 5149 2064 5155 2116
rect 5005 1904 5011 1916
rect 5053 1904 5059 1996
rect 5069 1984 5075 2036
rect 5133 1884 5139 1936
rect 5165 1903 5171 2116
rect 5245 2084 5251 2116
rect 5293 2084 5299 2276
rect 5197 1924 5203 2036
rect 5156 1897 5171 1903
rect 4733 1557 4755 1563
rect 4701 1544 4707 1556
rect 4669 1124 4675 1176
rect 4701 1084 4707 1316
rect 4717 1184 4723 1496
rect 4749 1364 4755 1557
rect 4797 1424 4803 1516
rect 4813 1184 4819 1356
rect 4829 1264 4835 1336
rect 4509 924 4515 1056
rect 4525 1044 4531 1056
rect 4621 984 4627 1056
rect 4685 944 4691 976
rect 4541 844 4547 876
rect 4605 864 4611 936
rect 4442 814 4454 816
rect 4427 806 4429 814
rect 4437 806 4439 814
rect 4447 806 4449 814
rect 4457 806 4459 814
rect 4467 806 4469 814
rect 4442 804 4454 806
rect 4093 364 4099 376
rect 4125 343 4131 396
rect 4221 384 4227 476
rect 4221 364 4227 376
rect 4109 337 4131 343
rect 4045 304 4051 316
rect 3965 264 3971 276
rect 4013 164 4019 196
rect 4029 184 4035 236
rect 3965 144 3971 156
rect 4045 144 4051 156
rect 3613 117 3628 123
rect 2317 84 2323 96
rect 3613 84 3619 117
rect 4061 104 4067 256
rect 4077 184 4083 276
rect 4077 144 4083 176
rect 4093 123 4099 216
rect 4084 117 4099 123
rect 4109 104 4115 337
rect 4157 284 4163 356
rect 4285 304 4291 516
rect 4317 504 4323 516
rect 4333 404 4339 656
rect 4381 484 4387 636
rect 4413 524 4419 756
rect 4493 604 4499 816
rect 4525 784 4531 836
rect 4701 804 4707 1056
rect 4749 904 4755 916
rect 4765 904 4771 1116
rect 4845 1104 4851 1496
rect 4893 1484 4899 1756
rect 4925 1644 4931 1756
rect 4941 1684 4947 1696
rect 4861 1304 4867 1356
rect 4893 1104 4899 1456
rect 4925 1383 4931 1536
rect 4957 1484 4963 1876
rect 5021 1784 5027 1876
rect 5069 1744 5075 1756
rect 4989 1724 4995 1736
rect 5133 1724 5139 1856
rect 4973 1604 4979 1636
rect 5197 1544 5203 1916
rect 4989 1424 4995 1496
rect 4909 1377 4931 1383
rect 4909 1364 4915 1377
rect 4909 1324 4915 1356
rect 4925 1344 4931 1356
rect 4989 1304 4995 1318
rect 4925 1084 4931 1196
rect 4724 897 4739 903
rect 4733 724 4739 897
rect 4637 702 4643 716
rect 4733 704 4739 716
rect 4637 544 4643 656
rect 4442 414 4454 416
rect 4427 406 4429 414
rect 4437 406 4439 414
rect 4447 406 4449 414
rect 4457 406 4459 414
rect 4467 406 4469 414
rect 4442 404 4454 406
rect 4125 124 4131 236
rect 4157 184 4163 256
rect 4173 224 4179 236
rect 4173 164 4179 196
rect 4253 124 4259 156
rect 4285 143 4291 296
rect 4333 264 4339 296
rect 4381 204 4387 256
rect 4381 164 4387 196
rect 4276 137 4291 143
rect 4493 124 4499 196
rect 4509 143 4515 436
rect 4589 244 4595 296
rect 4637 284 4643 536
rect 4653 526 4659 596
rect 4717 544 4723 576
rect 4685 464 4691 536
rect 4717 384 4723 516
rect 4733 503 4739 696
rect 4749 564 4755 656
rect 4733 497 4748 503
rect 4669 284 4675 376
rect 4765 303 4771 876
rect 4781 724 4787 1036
rect 4797 924 4803 936
rect 4797 864 4803 876
rect 4813 784 4819 856
rect 4797 704 4803 736
rect 4781 664 4787 676
rect 4813 624 4819 676
rect 4797 584 4803 596
rect 4781 504 4787 536
rect 4813 384 4819 516
rect 4829 504 4835 1056
rect 4845 924 4851 1076
rect 4893 1003 4899 1056
rect 4957 1023 4963 1094
rect 4877 997 4899 1003
rect 4941 1017 4963 1023
rect 4845 804 4851 896
rect 4861 784 4867 876
rect 4877 684 4883 997
rect 4941 984 4947 1017
rect 4893 944 4899 976
rect 4925 903 4931 956
rect 4909 897 4931 903
rect 4861 544 4867 616
rect 4877 583 4883 656
rect 4877 577 4899 583
rect 4829 364 4835 496
rect 4861 384 4867 516
rect 4765 297 4787 303
rect 4717 277 4732 283
rect 4717 244 4723 277
rect 4717 184 4723 236
rect 4557 144 4563 156
rect 4509 137 4531 143
rect 557 -17 563 36
rect 541 -23 563 -17
rect 701 -17 707 36
rect 1434 14 1446 16
rect 1419 6 1421 14
rect 1429 6 1431 14
rect 1439 6 1441 14
rect 1449 6 1451 14
rect 1459 6 1461 14
rect 1434 4 1446 6
rect 2205 -17 2211 36
rect 2493 -17 2499 36
rect 2541 -17 2547 36
rect 3085 -17 3091 36
rect 701 -23 723 -17
rect 2205 -23 2227 -17
rect 2493 -23 2515 -17
rect 2541 -23 2563 -17
rect 3069 -23 3091 -17
rect 3101 -17 3107 36
rect 3181 -17 3187 36
rect 3101 -23 3123 -17
rect 3165 -23 3187 -17
rect 3197 -17 3203 36
rect 3197 -23 3219 -17
rect 3501 -23 3507 16
rect 3565 -23 3571 16
rect 3661 -23 3667 16
rect 3709 -17 3715 36
rect 3693 -23 3715 -17
rect 3757 -23 3763 96
rect 3997 -23 4003 96
rect 4061 -23 4067 16
rect 4109 -23 4115 96
rect 4442 14 4454 16
rect 4427 6 4429 14
rect 4437 6 4439 14
rect 4447 6 4449 14
rect 4457 6 4459 14
rect 4467 6 4469 14
rect 4442 4 4454 6
rect 4525 -17 4531 137
rect 4685 124 4691 136
rect 4733 104 4739 256
rect 4749 144 4755 156
rect 4509 -23 4531 -17
rect 4589 -23 4595 96
rect 4733 -17 4739 96
rect 4717 -23 4739 -17
rect 4781 -23 4787 297
rect 4797 184 4803 216
rect 4813 184 4819 336
rect 4893 284 4899 577
rect 4909 564 4915 897
rect 4957 744 4963 936
rect 5005 804 5011 1516
rect 5101 1364 5107 1496
rect 5117 1484 5123 1516
rect 5165 1444 5171 1456
rect 5133 1424 5139 1436
rect 5021 944 5027 1136
rect 5053 1084 5059 1316
rect 5085 1184 5091 1316
rect 5197 1284 5203 1536
rect 5213 1524 5219 1916
rect 5229 1844 5235 1876
rect 5245 1804 5251 1856
rect 5245 1783 5251 1796
rect 5236 1777 5251 1783
rect 5245 1744 5251 1777
rect 5261 1724 5267 2076
rect 5277 1904 5283 1916
rect 5293 1724 5299 2036
rect 5309 1904 5315 2316
rect 5325 2304 5331 2416
rect 5373 2324 5379 2376
rect 5373 2304 5379 2316
rect 5325 2124 5331 2136
rect 5341 2124 5347 2296
rect 5357 2264 5363 2276
rect 5405 2264 5411 2396
rect 5325 1884 5331 2036
rect 5341 2024 5347 2116
rect 5373 1984 5379 2216
rect 5405 2124 5411 2136
rect 5421 2123 5427 2376
rect 5437 2323 5443 2336
rect 5469 2324 5475 2556
rect 5485 2424 5491 2637
rect 5501 2524 5507 2676
rect 5517 2604 5523 3036
rect 5597 2824 5603 3077
rect 5629 2984 5635 3036
rect 5645 2944 5651 2956
rect 5581 2664 5587 2736
rect 5501 2464 5507 2516
rect 5565 2504 5571 2516
rect 5581 2424 5587 2436
rect 5437 2317 5459 2323
rect 5453 2304 5459 2317
rect 5540 2317 5555 2323
rect 5437 2244 5443 2296
rect 5501 2284 5507 2296
rect 5460 2277 5475 2283
rect 5469 2263 5475 2277
rect 5533 2283 5539 2316
rect 5524 2277 5539 2283
rect 5469 2257 5500 2263
rect 5469 2184 5475 2236
rect 5485 2124 5491 2136
rect 5421 2117 5436 2123
rect 5389 1984 5395 2036
rect 5341 1904 5347 1976
rect 5213 1504 5219 1516
rect 5229 1504 5235 1556
rect 5245 1404 5251 1436
rect 5261 1424 5267 1716
rect 5293 1664 5299 1696
rect 5309 1663 5315 1736
rect 5389 1724 5395 1816
rect 5373 1703 5379 1716
rect 5373 1697 5395 1703
rect 5389 1684 5395 1697
rect 5405 1684 5411 2116
rect 5421 1884 5427 1996
rect 5300 1657 5315 1663
rect 5277 1504 5283 1576
rect 5421 1564 5427 1616
rect 5405 1524 5411 1556
rect 5293 1484 5299 1496
rect 5325 1484 5331 1496
rect 5213 1324 5219 1376
rect 5277 1364 5283 1476
rect 5069 944 5075 1176
rect 5101 1064 5107 1256
rect 5133 1144 5139 1236
rect 5181 1184 5187 1236
rect 5133 1104 5139 1116
rect 5117 984 5123 1016
rect 5101 924 5107 956
rect 5037 784 5043 896
rect 5133 884 5139 1056
rect 5213 1044 5219 1096
rect 5213 944 5219 956
rect 5229 924 5235 976
rect 5245 944 5251 1136
rect 5149 904 5155 916
rect 5181 884 5187 916
rect 5261 804 5267 1096
rect 5309 964 5315 1436
rect 5341 1323 5347 1436
rect 5332 1317 5347 1323
rect 5325 1084 5331 1136
rect 5389 1104 5395 1516
rect 5437 1503 5443 2116
rect 5485 2044 5491 2116
rect 5517 2104 5523 2116
rect 5453 1864 5459 1896
rect 5469 1884 5475 2036
rect 5533 1924 5539 2036
rect 5549 1964 5555 2317
rect 5581 2264 5587 2276
rect 5581 2124 5587 2156
rect 5565 2104 5571 2116
rect 5597 2064 5603 2456
rect 5613 2384 5619 2836
rect 5645 2824 5651 2936
rect 5709 2724 5715 3096
rect 5725 3084 5731 3116
rect 5725 2804 5731 3076
rect 5645 2684 5651 2694
rect 5709 2564 5715 2696
rect 5741 2604 5747 3137
rect 5757 3104 5763 3116
rect 5805 3104 5811 3476
rect 5837 3264 5843 3676
rect 5853 3584 5859 3896
rect 5949 3884 5955 4116
rect 5885 3744 5891 3836
rect 5901 3804 5907 3876
rect 5946 3814 5958 3816
rect 5931 3806 5933 3814
rect 5941 3806 5943 3814
rect 5951 3806 5953 3814
rect 5961 3806 5963 3814
rect 5971 3806 5973 3814
rect 5946 3804 5958 3806
rect 5997 3783 6003 4397
rect 6045 4264 6051 4296
rect 6013 4144 6019 4216
rect 6029 4184 6035 4256
rect 6029 4084 6035 4156
rect 6061 4124 6067 4496
rect 6077 4324 6083 4516
rect 6109 4424 6115 4556
rect 6125 4544 6131 4696
rect 6157 4684 6163 4696
rect 6173 4683 6179 4716
rect 6205 4704 6211 4836
rect 6333 4704 6339 4716
rect 6205 4684 6211 4696
rect 6164 4677 6179 4683
rect 6301 4664 6307 4696
rect 6141 4584 6147 4616
rect 6237 4584 6243 4616
rect 6196 4537 6243 4543
rect 6141 4524 6147 4536
rect 6237 4524 6243 4537
rect 6173 4464 6179 4516
rect 6253 4444 6259 4556
rect 6157 4384 6163 4416
rect 6093 4223 6099 4376
rect 6269 4324 6275 4576
rect 6285 4504 6291 4516
rect 6301 4344 6307 4496
rect 6173 4304 6179 4316
rect 6221 4264 6227 4276
rect 6093 4217 6115 4223
rect 6077 4144 6083 4156
rect 6045 4024 6051 4076
rect 6061 4024 6067 4116
rect 6045 3964 6051 3996
rect 6061 3984 6067 4016
rect 6029 3904 6035 3956
rect 6109 3944 6115 4217
rect 6205 4204 6211 4256
rect 6221 4224 6227 4236
rect 6221 4183 6227 4216
rect 6205 4177 6227 4183
rect 6205 4144 6211 4177
rect 6013 3824 6019 3856
rect 6029 3784 6035 3896
rect 6061 3804 6067 3916
rect 6077 3824 6083 3876
rect 6109 3864 6115 3916
rect 5981 3777 6003 3783
rect 5869 3724 5875 3736
rect 5885 3284 5891 3736
rect 5901 3424 5907 3496
rect 5965 3464 5971 3776
rect 5981 3604 5987 3777
rect 6093 3763 6099 3836
rect 6109 3784 6115 3856
rect 6093 3757 6115 3763
rect 6029 3664 6035 3696
rect 6045 3664 6051 3716
rect 6013 3584 6019 3596
rect 6061 3564 6067 3716
rect 6077 3684 6083 3716
rect 6061 3504 6067 3516
rect 5901 3383 5907 3416
rect 5946 3414 5958 3416
rect 5931 3406 5933 3414
rect 5941 3406 5943 3414
rect 5951 3406 5953 3414
rect 5961 3406 5963 3414
rect 5971 3406 5973 3414
rect 5946 3404 5958 3406
rect 5997 3384 6003 3496
rect 5901 3377 5916 3383
rect 5821 3124 5827 3156
rect 5885 3084 5891 3276
rect 6077 3264 6083 3656
rect 6093 3564 6099 3736
rect 6109 3703 6115 3757
rect 6125 3723 6131 3996
rect 6141 3924 6147 4136
rect 6221 4124 6227 4156
rect 6141 3804 6147 3896
rect 6173 3804 6179 4116
rect 6189 4064 6195 4116
rect 6221 4004 6227 4116
rect 6189 3904 6195 3956
rect 6221 3904 6227 3936
rect 6157 3724 6163 3776
rect 6125 3717 6147 3723
rect 6109 3697 6124 3703
rect 6093 3464 6099 3556
rect 6141 3503 6147 3717
rect 6173 3663 6179 3736
rect 6157 3657 6179 3663
rect 6157 3504 6163 3657
rect 6205 3644 6211 3896
rect 6221 3664 6227 3896
rect 6237 3864 6243 4316
rect 6269 4164 6275 4296
rect 6285 4144 6291 4276
rect 6317 4263 6323 4696
rect 6349 4683 6355 4716
rect 6381 4704 6387 4756
rect 6413 4724 6419 4856
rect 6340 4677 6355 4683
rect 6413 4683 6419 4716
rect 6429 4704 6435 4716
rect 6445 4704 6451 4916
rect 6541 4844 6547 4916
rect 6589 4724 6595 4736
rect 6404 4677 6419 4683
rect 6397 4544 6403 4656
rect 6413 4543 6419 4677
rect 6445 4624 6451 4696
rect 6477 4684 6483 4716
rect 6509 4684 6515 4696
rect 6621 4684 6627 4936
rect 6669 4924 6675 4936
rect 6685 4924 6691 4936
rect 6781 4924 6787 4936
rect 7005 4924 7011 5236
rect 7021 5023 7027 5316
rect 7085 5244 7091 5316
rect 7101 5304 7107 5316
rect 7277 5304 7283 5316
rect 7101 5044 7107 5296
rect 7117 5102 7123 5116
rect 7181 5064 7187 5136
rect 7197 5084 7203 5296
rect 7277 5104 7283 5216
rect 7213 5084 7219 5096
rect 7021 5017 7043 5023
rect 6765 4844 6771 4916
rect 6701 4764 6707 4836
rect 6797 4804 6803 4836
rect 6829 4784 6835 4916
rect 6861 4904 6867 4916
rect 6413 4537 6428 4543
rect 6333 4484 6339 4516
rect 6333 4304 6339 4476
rect 6349 4343 6355 4536
rect 6477 4524 6483 4616
rect 6365 4464 6371 4516
rect 6493 4344 6499 4536
rect 6509 4424 6515 4676
rect 6589 4524 6595 4616
rect 6525 4464 6531 4516
rect 6621 4464 6627 4516
rect 6349 4337 6364 4343
rect 6333 4284 6339 4296
rect 6557 4284 6563 4336
rect 6637 4304 6643 4316
rect 6653 4303 6659 4736
rect 6701 4664 6707 4696
rect 6669 4524 6675 4636
rect 6781 4624 6787 4636
rect 6749 4564 6755 4616
rect 6813 4584 6819 4696
rect 6861 4564 6867 4776
rect 6941 4684 6947 4696
rect 6925 4584 6931 4616
rect 7021 4584 7027 4596
rect 6701 4524 6707 4556
rect 6749 4524 6755 4536
rect 6829 4524 6835 4536
rect 6941 4524 6947 4536
rect 6957 4524 6963 4536
rect 6685 4484 6691 4516
rect 6717 4324 6723 4336
rect 6797 4304 6803 4316
rect 6653 4297 6668 4303
rect 6589 4284 6595 4296
rect 6317 4257 6339 4263
rect 6301 4164 6307 4196
rect 6269 4024 6275 4116
rect 6253 3984 6259 3996
rect 6253 3924 6259 3976
rect 6269 3884 6275 3956
rect 6285 3924 6291 4136
rect 6333 4123 6339 4257
rect 6349 4224 6355 4276
rect 6349 4144 6355 4176
rect 6365 4124 6371 4176
rect 6445 4144 6451 4216
rect 6388 4137 6403 4143
rect 6333 4117 6355 4123
rect 6301 3984 6307 4076
rect 6292 3897 6307 3903
rect 6301 3864 6307 3897
rect 6253 3764 6259 3776
rect 6125 3497 6147 3503
rect 6125 3464 6131 3497
rect 6093 3324 6099 3376
rect 6061 3257 6076 3263
rect 5789 3024 5795 3036
rect 5853 2984 5859 3036
rect 5869 2964 5875 3016
rect 5946 3014 5958 3016
rect 5931 3006 5933 3014
rect 5941 3006 5943 3014
rect 5951 3006 5953 3014
rect 5961 3006 5963 3014
rect 5971 3006 5973 3014
rect 5946 3004 5958 3006
rect 5821 2924 5827 2936
rect 5821 2904 5827 2916
rect 5757 2704 5763 2836
rect 5789 2764 5795 2836
rect 5693 2524 5699 2556
rect 5613 2304 5619 2316
rect 5661 2304 5667 2316
rect 5677 2284 5683 2296
rect 5693 2264 5699 2336
rect 5709 2284 5715 2556
rect 5773 2484 5779 2716
rect 5789 2624 5795 2716
rect 5805 2704 5811 2756
rect 5821 2664 5827 2796
rect 5805 2524 5811 2596
rect 5821 2524 5827 2616
rect 5805 2464 5811 2516
rect 5725 2264 5731 2296
rect 5773 2284 5779 2416
rect 5796 2317 5811 2323
rect 5805 2304 5811 2317
rect 5629 2184 5635 2236
rect 5741 2224 5747 2276
rect 5773 2264 5779 2276
rect 5613 2144 5619 2156
rect 5661 2144 5667 2156
rect 5597 1903 5603 2056
rect 5588 1897 5603 1903
rect 5485 1664 5491 1736
rect 5517 1724 5523 1896
rect 5549 1864 5555 1896
rect 5549 1843 5555 1856
rect 5540 1837 5555 1843
rect 5501 1664 5507 1716
rect 5549 1643 5555 1756
rect 5565 1724 5571 1876
rect 5581 1864 5587 1876
rect 5613 1863 5619 2136
rect 5677 2124 5683 2196
rect 5741 2164 5747 2216
rect 5645 1944 5651 2116
rect 5645 1904 5651 1936
rect 5661 1903 5667 2016
rect 5741 2004 5747 2156
rect 5757 2124 5763 2176
rect 5773 2164 5779 2256
rect 5709 1924 5715 1956
rect 5661 1897 5676 1903
rect 5645 1863 5651 1876
rect 5613 1857 5651 1863
rect 5645 1784 5651 1857
rect 5581 1744 5587 1756
rect 5597 1724 5603 1776
rect 5661 1744 5667 1796
rect 5629 1737 5644 1743
rect 5629 1704 5635 1737
rect 5677 1724 5683 1896
rect 5709 1764 5715 1916
rect 5773 1904 5779 2076
rect 5789 2064 5795 2296
rect 5821 2264 5827 2516
rect 5837 2424 5843 2916
rect 5885 2884 5891 2916
rect 5901 2904 5907 2996
rect 5981 2904 5987 2936
rect 5885 2704 5891 2876
rect 5933 2784 5939 2796
rect 5901 2704 5907 2736
rect 5997 2704 6003 3216
rect 6045 3104 6051 3236
rect 6061 3063 6067 3257
rect 6045 3057 6067 3063
rect 6029 2903 6035 2916
rect 6013 2897 6035 2903
rect 6013 2804 6019 2897
rect 6029 2764 6035 2836
rect 5853 2644 5859 2696
rect 5869 2684 5875 2696
rect 5869 2584 5875 2656
rect 5946 2614 5958 2616
rect 5931 2606 5933 2614
rect 5941 2606 5943 2614
rect 5951 2606 5953 2614
rect 5961 2606 5963 2614
rect 5971 2606 5973 2614
rect 5946 2604 5958 2606
rect 5837 2204 5843 2336
rect 5869 2224 5875 2296
rect 5885 2184 5891 2376
rect 5869 2144 5875 2176
rect 5885 2104 5891 2176
rect 5901 2084 5907 2516
rect 5981 2504 5987 2516
rect 5917 2284 5923 2296
rect 5946 2214 5958 2216
rect 5931 2206 5933 2214
rect 5941 2206 5943 2214
rect 5951 2206 5953 2214
rect 5961 2206 5963 2214
rect 5971 2206 5973 2214
rect 5946 2204 5958 2206
rect 5789 1904 5795 1976
rect 5757 1864 5763 1896
rect 5725 1844 5731 1856
rect 5725 1764 5731 1836
rect 5757 1824 5763 1836
rect 5773 1824 5779 1896
rect 5837 1883 5843 1936
rect 5853 1904 5859 1936
rect 5885 1904 5891 1916
rect 5933 1884 5939 1956
rect 5837 1877 5852 1883
rect 5645 1644 5651 1716
rect 5709 1704 5715 1756
rect 5757 1724 5763 1816
rect 5805 1723 5811 1836
rect 5821 1724 5827 1756
rect 5853 1744 5859 1776
rect 5869 1724 5875 1816
rect 5901 1784 5907 1876
rect 5965 1864 5971 2176
rect 5981 2124 5987 2136
rect 5981 1864 5987 2116
rect 5946 1814 5958 1816
rect 5931 1806 5933 1814
rect 5941 1806 5943 1814
rect 5951 1806 5953 1814
rect 5961 1806 5963 1814
rect 5971 1806 5973 1814
rect 5946 1804 5958 1806
rect 5796 1717 5811 1723
rect 5876 1717 5891 1723
rect 5693 1664 5699 1696
rect 5533 1637 5555 1643
rect 5517 1504 5523 1596
rect 5533 1504 5539 1637
rect 5597 1524 5603 1636
rect 5757 1543 5763 1716
rect 5741 1537 5763 1543
rect 5428 1497 5443 1503
rect 5533 1484 5539 1496
rect 5517 1463 5523 1476
rect 5517 1457 5564 1463
rect 5405 1384 5411 1456
rect 5421 1324 5427 1416
rect 5437 1324 5443 1436
rect 5453 1404 5459 1436
rect 5501 1424 5507 1456
rect 5501 1324 5507 1416
rect 5533 1404 5539 1436
rect 5581 1424 5587 1436
rect 5533 1324 5539 1396
rect 5581 1324 5587 1416
rect 5645 1364 5651 1496
rect 5693 1484 5699 1496
rect 5693 1324 5699 1416
rect 5405 1124 5411 1236
rect 5453 1104 5459 1176
rect 5469 1164 5475 1236
rect 5517 1184 5523 1316
rect 5533 1184 5539 1196
rect 5565 1184 5571 1236
rect 5629 1184 5635 1316
rect 5661 1244 5667 1316
rect 5693 1304 5699 1316
rect 5396 1097 5404 1103
rect 5357 1084 5363 1096
rect 5405 1044 5411 1096
rect 5437 1064 5443 1076
rect 5309 944 5315 956
rect 5389 924 5395 996
rect 5421 964 5427 1056
rect 5453 964 5459 1076
rect 5469 944 5475 956
rect 5485 944 5491 1116
rect 5517 1103 5523 1176
rect 5517 1097 5532 1103
rect 5533 1064 5539 1096
rect 5581 1084 5587 1116
rect 5597 1104 5603 1176
rect 5501 964 5507 1036
rect 5453 924 5459 936
rect 5517 924 5523 1016
rect 5533 944 5539 956
rect 5549 944 5555 976
rect 5581 964 5587 1076
rect 5629 1063 5635 1096
rect 5645 1084 5651 1196
rect 5677 1104 5683 1176
rect 5661 1084 5667 1096
rect 5693 1084 5699 1296
rect 5709 1124 5715 1256
rect 5725 1184 5731 1396
rect 5741 1204 5747 1537
rect 5805 1504 5811 1616
rect 5869 1504 5875 1596
rect 5885 1584 5891 1717
rect 5901 1704 5907 1756
rect 5997 1743 6003 2696
rect 6013 2524 6019 2536
rect 6029 2524 6035 2536
rect 6029 2363 6035 2476
rect 6045 2384 6051 3057
rect 6093 3044 6099 3056
rect 6061 2924 6067 3036
rect 6077 2944 6083 3016
rect 6109 2984 6115 3456
rect 6141 3443 6147 3476
rect 6157 3444 6163 3496
rect 6125 3437 6147 3443
rect 6125 3344 6131 3437
rect 6189 3384 6195 3636
rect 6221 3524 6227 3636
rect 6189 3364 6195 3376
rect 6125 3084 6131 3336
rect 6157 3324 6163 3336
rect 6189 3104 6195 3256
rect 6093 2784 6099 2956
rect 6109 2704 6115 2736
rect 6125 2704 6131 3036
rect 6141 2864 6147 3096
rect 6157 2884 6163 2936
rect 6173 2924 6179 3076
rect 6173 2703 6179 2916
rect 6157 2697 6179 2703
rect 6189 2703 6195 2976
rect 6221 2924 6227 3456
rect 6253 3424 6259 3756
rect 6285 3744 6291 3856
rect 6285 3504 6291 3736
rect 6317 3724 6323 4016
rect 6349 3904 6355 4117
rect 6397 4104 6403 4137
rect 6397 4004 6403 4096
rect 6429 4064 6435 4116
rect 6461 4044 6467 4136
rect 6477 4104 6483 4116
rect 6301 3684 6307 3716
rect 6333 3664 6339 3896
rect 6349 3784 6355 3896
rect 6365 3884 6371 3916
rect 6381 3764 6387 3896
rect 6397 3744 6403 3996
rect 6413 3904 6419 3936
rect 6413 3784 6419 3816
rect 6461 3784 6467 4036
rect 6477 4004 6483 4096
rect 6493 3904 6499 4276
rect 6525 4264 6531 4276
rect 6509 4084 6515 4196
rect 6573 4144 6579 4196
rect 6548 4117 6556 4123
rect 6541 3924 6547 4116
rect 6573 4024 6579 4136
rect 6621 3984 6627 4276
rect 6653 4144 6659 4256
rect 6509 3904 6515 3916
rect 6573 3904 6579 3936
rect 6653 3904 6659 4076
rect 6669 3984 6675 4296
rect 6845 4284 6851 4516
rect 6957 4284 6963 4516
rect 6717 4244 6723 4276
rect 6829 4204 6835 4276
rect 6701 4104 6707 4116
rect 6781 4084 6787 4116
rect 6797 4104 6803 4116
rect 6493 3784 6499 3856
rect 6509 3723 6515 3896
rect 6621 3884 6627 3896
rect 6557 3764 6563 3816
rect 6573 3804 6579 3876
rect 6637 3844 6643 3896
rect 6669 3884 6675 3896
rect 6749 3884 6755 3936
rect 6781 3904 6787 3916
rect 6509 3717 6531 3723
rect 6429 3704 6435 3716
rect 6349 3564 6355 3676
rect 6493 3604 6499 3716
rect 6397 3504 6403 3556
rect 6413 3504 6419 3536
rect 6285 3344 6291 3496
rect 6317 3326 6323 3396
rect 6349 3324 6355 3336
rect 6244 3137 6259 3143
rect 6237 3104 6243 3116
rect 6253 3104 6259 3137
rect 6397 3104 6403 3496
rect 6445 3384 6451 3396
rect 6413 3324 6419 3336
rect 6445 3184 6451 3256
rect 6461 3164 6467 3336
rect 6477 3324 6483 3416
rect 6525 3384 6531 3717
rect 6541 3704 6547 3736
rect 6605 3684 6611 3736
rect 6621 3724 6627 3836
rect 6701 3764 6707 3856
rect 6653 3704 6659 3736
rect 6701 3684 6707 3756
rect 6717 3744 6723 3776
rect 6733 3724 6739 3836
rect 6781 3624 6787 3896
rect 6813 3724 6819 3916
rect 6845 3884 6851 4276
rect 6877 4124 6883 4236
rect 6925 4224 6931 4276
rect 6925 4184 6931 4216
rect 6893 4024 6899 4116
rect 6941 4104 6947 4116
rect 6941 4084 6947 4096
rect 6845 3764 6851 3876
rect 6845 3717 6860 3723
rect 6829 3624 6835 3716
rect 6717 3584 6723 3616
rect 6637 3524 6643 3536
rect 6541 3502 6547 3516
rect 6605 3484 6611 3496
rect 6653 3484 6659 3516
rect 6685 3504 6691 3536
rect 6845 3503 6851 3717
rect 6877 3704 6883 3716
rect 6877 3564 6883 3696
rect 6845 3497 6867 3503
rect 6493 3324 6499 3376
rect 6541 3324 6547 3336
rect 6573 3324 6579 3476
rect 6477 3284 6483 3316
rect 6493 3264 6499 3316
rect 6525 3124 6531 3236
rect 6573 3184 6579 3236
rect 6573 3124 6579 3176
rect 6477 3104 6483 3116
rect 6269 3083 6275 3096
rect 6301 3084 6307 3096
rect 6333 3084 6339 3096
rect 6260 3077 6275 3083
rect 6285 2924 6291 3076
rect 6317 3064 6323 3076
rect 6365 3044 6371 3096
rect 6525 3084 6531 3096
rect 6301 2984 6307 2996
rect 6333 2924 6339 2996
rect 6365 2984 6371 3016
rect 6381 2964 6387 3076
rect 6413 2944 6419 2956
rect 6429 2923 6435 3076
rect 6461 3044 6467 3076
rect 6493 3057 6508 3063
rect 6477 2944 6483 3036
rect 6413 2917 6435 2923
rect 6205 2884 6211 2896
rect 6189 2697 6204 2703
rect 6061 2624 6067 2696
rect 6125 2684 6131 2696
rect 6061 2564 6067 2616
rect 6125 2564 6131 2596
rect 6141 2584 6147 2616
rect 6125 2524 6131 2556
rect 6093 2484 6099 2516
rect 6029 2357 6051 2363
rect 6029 2164 6035 2276
rect 6045 2184 6051 2357
rect 6061 2224 6067 2256
rect 6061 2184 6067 2216
rect 6045 2004 6051 2096
rect 6013 1904 6019 1916
rect 6029 1904 6035 1976
rect 6045 1864 6051 1896
rect 6061 1744 6067 2076
rect 6077 2024 6083 2376
rect 6109 2304 6115 2316
rect 6141 2204 6147 2456
rect 6157 2324 6163 2697
rect 6093 2044 6099 2116
rect 6077 1924 6083 2016
rect 6109 2004 6115 2136
rect 6125 2083 6131 2136
rect 6125 2077 6147 2083
rect 6125 1984 6131 2036
rect 6093 1944 6099 1976
rect 6077 1824 6083 1916
rect 6093 1904 6099 1936
rect 5981 1737 6003 1743
rect 5901 1564 5907 1596
rect 5981 1524 5987 1737
rect 5997 1664 6003 1716
rect 6045 1644 6051 1716
rect 5997 1544 6003 1616
rect 5805 1484 5811 1496
rect 5773 1384 5779 1456
rect 5773 1324 5779 1356
rect 5789 1324 5795 1376
rect 5725 1104 5731 1136
rect 5773 1084 5779 1116
rect 5789 1104 5795 1156
rect 5709 1077 5724 1083
rect 5709 1063 5715 1077
rect 5741 1077 5756 1083
rect 5629 1057 5715 1063
rect 5677 984 5683 1016
rect 5197 784 5203 796
rect 5117 724 5123 776
rect 5309 764 5315 916
rect 5341 904 5347 916
rect 4909 484 4915 516
rect 4941 444 4947 616
rect 4957 504 4963 696
rect 5021 544 5027 656
rect 5117 624 5123 716
rect 5149 664 5155 676
rect 5261 664 5267 676
rect 5181 564 5187 656
rect 5213 604 5219 656
rect 5229 564 5235 656
rect 5293 624 5299 716
rect 5325 684 5331 736
rect 5117 544 5123 556
rect 5373 544 5379 616
rect 5405 604 5411 916
rect 5469 903 5475 916
rect 5453 897 5475 903
rect 5453 884 5459 897
rect 5453 704 5459 796
rect 5501 704 5507 916
rect 5517 784 5523 896
rect 5533 784 5539 936
rect 5565 924 5571 936
rect 5661 924 5667 936
rect 5725 924 5731 1056
rect 5741 984 5747 1077
rect 5757 1064 5763 1076
rect 5533 744 5539 776
rect 5549 764 5555 796
rect 5453 684 5459 696
rect 5485 544 5491 576
rect 4957 364 4963 476
rect 5021 464 5027 536
rect 4973 384 4979 436
rect 5021 384 5027 456
rect 4797 144 4803 176
rect 4829 123 4835 256
rect 4845 204 4851 256
rect 4861 183 4867 196
rect 4909 184 4915 236
rect 4925 184 4931 236
rect 4852 177 4867 183
rect 4813 117 4835 123
rect 4813 103 4819 117
rect 4804 97 4819 103
rect 4813 -23 4819 97
rect 4829 84 4835 96
rect 4861 -23 4867 76
rect 4893 -23 4899 36
rect 4941 -17 4947 356
rect 4957 304 4963 356
rect 4925 -23 4947 -17
rect 4957 -23 4963 236
rect 4973 126 4979 256
rect 4989 244 4995 256
rect 5069 183 5075 276
rect 5117 184 5123 476
rect 5181 344 5187 536
rect 5213 504 5219 536
rect 5245 517 5260 523
rect 5149 324 5155 336
rect 5069 177 5107 183
rect 5069 144 5075 177
rect 5037 124 5043 136
rect 5053 97 5068 103
rect 5053 -23 5059 97
rect 5101 -23 5107 177
rect 5117 124 5123 136
rect 5117 104 5123 116
rect 5149 103 5155 236
rect 5165 184 5171 296
rect 5197 224 5203 276
rect 5213 184 5219 456
rect 5245 384 5251 517
rect 5277 364 5283 516
rect 5373 504 5379 536
rect 5181 124 5187 136
rect 5229 124 5235 236
rect 5245 144 5251 336
rect 5277 304 5283 356
rect 5389 304 5395 516
rect 5437 484 5443 536
rect 5501 384 5507 696
rect 5421 323 5427 336
rect 5421 317 5436 323
rect 5309 224 5315 236
rect 5277 164 5283 216
rect 5357 184 5363 276
rect 5373 264 5379 296
rect 5549 284 5555 756
rect 5565 704 5571 896
rect 5613 724 5619 916
rect 5629 804 5635 916
rect 5581 624 5587 636
rect 5645 544 5651 676
rect 5709 624 5715 694
rect 5741 664 5747 676
rect 5773 644 5779 696
rect 5677 564 5683 616
rect 5741 584 5747 616
rect 5469 204 5475 276
rect 5485 183 5491 256
rect 5476 177 5491 183
rect 5549 124 5555 136
rect 5581 124 5587 536
rect 5773 524 5779 616
rect 5805 543 5811 1476
rect 5869 1444 5875 1496
rect 5837 1326 5843 1436
rect 5885 1404 5891 1436
rect 5901 1344 5907 1516
rect 5917 1504 5923 1516
rect 5981 1443 5987 1516
rect 5997 1504 6003 1536
rect 5981 1437 6003 1443
rect 5946 1414 5958 1416
rect 5931 1406 5933 1414
rect 5941 1406 5943 1414
rect 5951 1406 5953 1414
rect 5961 1406 5963 1414
rect 5971 1406 5973 1414
rect 5946 1404 5958 1406
rect 5837 1084 5843 1096
rect 5853 1064 5859 1076
rect 5837 704 5843 1036
rect 5869 963 5875 1156
rect 5885 1104 5891 1196
rect 5853 957 5875 963
rect 5853 924 5859 957
rect 5837 684 5843 696
rect 5869 684 5875 936
rect 5901 924 5907 1336
rect 5949 1304 5955 1356
rect 5917 1124 5923 1236
rect 5981 1104 5987 1176
rect 5946 1014 5958 1016
rect 5931 1006 5933 1014
rect 5941 1006 5943 1014
rect 5951 1006 5953 1014
rect 5961 1006 5963 1014
rect 5971 1006 5973 1014
rect 5946 1004 5958 1006
rect 5997 943 6003 1437
rect 6013 1344 6019 1636
rect 6061 1564 6067 1716
rect 6077 1624 6083 1776
rect 6093 1724 6099 1796
rect 6125 1764 6131 1936
rect 6141 1924 6147 2077
rect 6157 1964 6163 2276
rect 6173 2264 6179 2296
rect 6173 2184 6179 2196
rect 6173 2104 6179 2176
rect 6205 2164 6211 2516
rect 6221 2304 6227 2916
rect 6269 2723 6275 2736
rect 6253 2717 6275 2723
rect 6253 2704 6259 2717
rect 6253 2644 6259 2676
rect 6253 2484 6259 2516
rect 6269 2304 6275 2696
rect 6301 2664 6307 2776
rect 6317 2724 6323 2896
rect 6317 2684 6323 2716
rect 6333 2564 6339 2776
rect 6365 2704 6371 2876
rect 6381 2684 6387 2896
rect 6397 2884 6403 2916
rect 6397 2704 6403 2736
rect 6365 2644 6371 2676
rect 6413 2643 6419 2917
rect 6429 2684 6435 2696
rect 6445 2684 6451 2916
rect 6461 2884 6467 2916
rect 6493 2664 6499 3057
rect 6541 3004 6547 3116
rect 6557 2943 6563 3076
rect 6573 3024 6579 3096
rect 6605 3084 6611 3096
rect 6637 3084 6643 3096
rect 6589 3064 6595 3076
rect 6557 2937 6579 2943
rect 6573 2924 6579 2937
rect 6509 2864 6515 2916
rect 6525 2684 6531 2696
rect 6413 2637 6435 2643
rect 6413 2584 6419 2616
rect 6301 2544 6307 2556
rect 6429 2524 6435 2637
rect 6509 2624 6515 2676
rect 6541 2603 6547 2836
rect 6557 2664 6563 2716
rect 6525 2597 6547 2603
rect 6237 2284 6243 2296
rect 6237 2224 6243 2256
rect 6269 2184 6275 2296
rect 6205 2144 6211 2156
rect 6173 1863 6179 2076
rect 6237 1924 6243 1996
rect 6173 1857 6195 1863
rect 6173 1724 6179 1736
rect 6141 1644 6147 1716
rect 6109 1604 6115 1636
rect 6029 1444 6035 1536
rect 6045 1504 6051 1516
rect 6093 1504 6099 1556
rect 6141 1504 6147 1516
rect 6125 1484 6131 1496
rect 6029 1344 6035 1436
rect 6077 1424 6083 1436
rect 6061 1344 6067 1356
rect 6045 1324 6051 1336
rect 6013 1184 6019 1216
rect 6029 1104 6035 1296
rect 6045 1104 6051 1256
rect 6061 1184 6067 1276
rect 6077 1204 6083 1276
rect 6093 1224 6099 1336
rect 6109 1324 6115 1396
rect 5997 937 6019 943
rect 5869 664 5875 676
rect 5796 537 5811 543
rect 5789 524 5795 536
rect 5821 524 5827 536
rect 5613 284 5619 476
rect 5789 344 5795 516
rect 5805 504 5811 516
rect 5748 297 5772 303
rect 5645 204 5651 296
rect 5821 284 5827 476
rect 5853 323 5859 496
rect 5844 317 5859 323
rect 5869 284 5875 576
rect 5885 324 5891 636
rect 5901 604 5907 896
rect 5981 864 5987 936
rect 5997 804 6003 916
rect 6013 804 6019 937
rect 5933 664 5939 676
rect 5997 664 6003 796
rect 6013 704 6019 756
rect 5946 614 5958 616
rect 5931 606 5933 614
rect 5941 606 5943 614
rect 5951 606 5953 614
rect 5961 606 5963 614
rect 5971 606 5973 614
rect 5946 604 5958 606
rect 5901 384 5907 596
rect 6013 564 6019 676
rect 6029 564 6035 1036
rect 6045 1024 6051 1096
rect 6077 1024 6083 1196
rect 6093 1124 6099 1176
rect 6093 1084 6099 1116
rect 6109 1044 6115 1276
rect 6141 1183 6147 1436
rect 6157 1304 6163 1716
rect 6189 1564 6195 1857
rect 6253 1783 6259 2136
rect 6301 2024 6307 2316
rect 6317 2304 6323 2376
rect 6381 2324 6387 2516
rect 6429 2504 6435 2516
rect 6445 2504 6451 2576
rect 6477 2557 6515 2563
rect 6477 2544 6483 2557
rect 6509 2544 6515 2557
rect 6493 2524 6499 2536
rect 6525 2524 6531 2597
rect 6541 2544 6547 2576
rect 6413 2403 6419 2436
rect 6413 2397 6435 2403
rect 6413 2304 6419 2376
rect 6333 2284 6339 2296
rect 6365 2264 6371 2296
rect 6381 2264 6387 2276
rect 6269 1917 6323 1923
rect 6269 1904 6275 1917
rect 6317 1904 6323 1917
rect 6253 1777 6268 1783
rect 6221 1744 6227 1756
rect 6221 1724 6227 1736
rect 6253 1704 6259 1736
rect 6269 1704 6275 1716
rect 6285 1684 6291 1796
rect 6301 1744 6307 1836
rect 6333 1804 6339 2016
rect 6381 1984 6387 2156
rect 6413 2144 6419 2176
rect 6429 2124 6435 2397
rect 6445 2304 6451 2456
rect 6541 2444 6547 2536
rect 6573 2523 6579 2916
rect 6589 2584 6595 3056
rect 6653 3044 6659 3076
rect 6669 3064 6675 3236
rect 6685 3144 6691 3496
rect 6701 3444 6707 3476
rect 6717 3184 6723 3318
rect 6749 3243 6755 3496
rect 6813 3484 6819 3496
rect 6765 3384 6771 3456
rect 6781 3364 6787 3436
rect 6813 3344 6819 3476
rect 6797 3304 6803 3316
rect 6733 3237 6755 3243
rect 6669 2943 6675 3056
rect 6653 2937 6675 2943
rect 6605 2864 6611 2916
rect 6621 2684 6627 2936
rect 6653 2924 6659 2937
rect 6669 2884 6675 2916
rect 6685 2763 6691 3136
rect 6701 3104 6707 3116
rect 6701 2924 6707 2996
rect 6733 2904 6739 3237
rect 6749 3084 6755 3116
rect 6669 2757 6691 2763
rect 6669 2724 6675 2757
rect 6621 2604 6627 2676
rect 6637 2644 6643 2676
rect 6685 2664 6691 2736
rect 6637 2583 6643 2636
rect 6628 2577 6643 2583
rect 6573 2517 6588 2523
rect 6653 2504 6659 2636
rect 6685 2524 6691 2556
rect 6461 2404 6467 2436
rect 6445 2284 6451 2296
rect 6445 2137 6460 2143
rect 6445 2124 6451 2137
rect 6461 2104 6467 2116
rect 6429 2004 6435 2076
rect 6429 1923 6435 1996
rect 6477 1944 6483 2416
rect 6509 2317 6524 2323
rect 6493 1944 6499 2316
rect 6509 2244 6515 2317
rect 6525 2244 6531 2296
rect 6541 2143 6547 2336
rect 6557 2324 6563 2496
rect 6701 2424 6707 2896
rect 6717 2744 6723 2836
rect 6749 2644 6755 3076
rect 6765 2844 6771 3096
rect 6781 2984 6787 3096
rect 6813 3064 6819 3336
rect 6829 3264 6835 3316
rect 6845 3104 6851 3236
rect 6861 3104 6867 3497
rect 6877 3464 6883 3556
rect 6893 3544 6899 3876
rect 6925 3744 6931 4036
rect 6941 3864 6947 4076
rect 6957 3844 6963 4116
rect 7005 3983 7011 4516
rect 7037 4104 7043 5017
rect 7053 4944 7059 4956
rect 7101 4944 7107 4956
rect 7101 4917 7116 4923
rect 7069 4604 7075 4836
rect 7085 4624 7091 4696
rect 7101 4544 7107 4917
rect 7149 4744 7155 4836
rect 7133 4684 7139 4696
rect 7133 4544 7139 4676
rect 7165 4663 7171 4936
rect 7165 4657 7187 4663
rect 7165 4604 7171 4636
rect 7101 4284 7107 4516
rect 7133 4303 7139 4516
rect 7149 4504 7155 4518
rect 7181 4464 7187 4657
rect 7197 4623 7203 5076
rect 7213 4964 7219 5076
rect 7357 5023 7363 5116
rect 7341 5017 7363 5023
rect 7245 4703 7251 4916
rect 7341 4883 7347 5017
rect 7341 4877 7363 4883
rect 7236 4697 7251 4703
rect 7197 4617 7219 4623
rect 7213 4544 7219 4617
rect 7181 4383 7187 4456
rect 7181 4377 7196 4383
rect 7133 4297 7148 4303
rect 7149 4284 7155 4296
rect 7053 4144 7059 4276
rect 7053 4124 7059 4136
rect 6989 3977 7011 3983
rect 6973 3904 6979 3916
rect 6925 3664 6931 3716
rect 6909 3504 6915 3636
rect 6909 3444 6915 3496
rect 6877 3124 6883 3136
rect 6813 3024 6819 3036
rect 6845 3004 6851 3096
rect 6861 3084 6867 3096
rect 6765 2604 6771 2836
rect 6797 2704 6803 2716
rect 6845 2684 6851 2916
rect 6877 2704 6883 3076
rect 6909 3044 6915 3076
rect 6925 3023 6931 3536
rect 6909 3017 6931 3023
rect 6893 2924 6899 2956
rect 6909 2884 6915 3017
rect 6925 2744 6931 2776
rect 6893 2704 6899 2736
rect 6893 2684 6899 2696
rect 6845 2664 6851 2676
rect 6877 2624 6883 2676
rect 6557 2284 6563 2296
rect 6573 2284 6579 2316
rect 6621 2304 6627 2396
rect 6701 2384 6707 2396
rect 6701 2304 6707 2376
rect 6589 2224 6595 2256
rect 6621 2204 6627 2296
rect 6653 2264 6659 2296
rect 6669 2264 6675 2276
rect 6685 2204 6691 2296
rect 6532 2137 6547 2143
rect 6429 1917 6444 1923
rect 6349 1864 6355 1876
rect 6397 1864 6403 1876
rect 6365 1764 6371 1856
rect 6429 1844 6435 1896
rect 6493 1884 6499 1916
rect 6493 1863 6499 1876
rect 6525 1864 6531 2136
rect 6541 1984 6547 1996
rect 6557 1884 6563 2176
rect 6685 2164 6691 2196
rect 6589 2124 6595 2136
rect 6621 2124 6627 2136
rect 6637 2124 6643 2156
rect 6717 2144 6723 2236
rect 6733 2204 6739 2236
rect 6573 2104 6579 2116
rect 6717 2104 6723 2116
rect 6669 1984 6675 2036
rect 6612 1937 6627 1943
rect 6605 1924 6611 1936
rect 6573 1884 6579 1896
rect 6477 1857 6499 1863
rect 6381 1724 6387 1816
rect 6429 1744 6435 1816
rect 6477 1724 6483 1857
rect 6493 1744 6499 1756
rect 6509 1724 6515 1856
rect 6557 1824 6563 1876
rect 6589 1723 6595 1796
rect 6605 1744 6611 1836
rect 6621 1744 6627 1937
rect 6685 1904 6691 2076
rect 6733 1904 6739 1916
rect 6749 1824 6755 2576
rect 6861 2544 6867 2596
rect 6877 2544 6883 2576
rect 6845 2504 6851 2516
rect 6845 2383 6851 2496
rect 6861 2384 6867 2536
rect 6877 2464 6883 2536
rect 6829 2377 6851 2383
rect 6797 2144 6803 2256
rect 6765 2104 6771 2136
rect 6781 2124 6787 2136
rect 6813 2124 6819 2296
rect 6829 2124 6835 2377
rect 6845 2244 6851 2296
rect 6781 2064 6787 2116
rect 6653 1784 6659 1796
rect 6669 1724 6675 1816
rect 6580 1717 6595 1723
rect 6237 1584 6243 1636
rect 6205 1464 6211 1496
rect 6221 1423 6227 1556
rect 6269 1523 6275 1536
rect 6285 1524 6291 1636
rect 6253 1517 6275 1523
rect 6253 1504 6259 1517
rect 6237 1477 6252 1483
rect 6237 1424 6243 1477
rect 6269 1464 6275 1496
rect 6301 1464 6307 1676
rect 6317 1484 6323 1656
rect 6349 1544 6355 1716
rect 6445 1704 6451 1716
rect 6493 1703 6499 1716
rect 6493 1697 6515 1703
rect 6365 1484 6371 1516
rect 6397 1504 6403 1516
rect 6413 1484 6419 1696
rect 6509 1684 6515 1697
rect 6477 1504 6483 1556
rect 6493 1504 6499 1636
rect 6573 1624 6579 1636
rect 6589 1624 6595 1696
rect 6605 1584 6611 1716
rect 6445 1484 6451 1496
rect 6253 1443 6259 1456
rect 6317 1443 6323 1456
rect 6253 1437 6323 1443
rect 6349 1424 6355 1476
rect 6212 1417 6227 1423
rect 6173 1324 6179 1356
rect 6205 1324 6211 1416
rect 6333 1344 6339 1376
rect 6173 1224 6179 1296
rect 6221 1244 6227 1336
rect 6349 1324 6355 1376
rect 6365 1344 6371 1476
rect 6381 1464 6387 1476
rect 6461 1464 6467 1496
rect 6493 1484 6499 1496
rect 6397 1397 6499 1403
rect 6397 1384 6403 1397
rect 6493 1384 6499 1397
rect 6413 1364 6419 1376
rect 6461 1364 6467 1376
rect 6397 1343 6403 1356
rect 6397 1337 6412 1343
rect 6141 1177 6163 1183
rect 6157 1164 6163 1177
rect 6141 1084 6147 1096
rect 6157 1084 6163 1156
rect 6141 1044 6147 1076
rect 6189 1063 6195 1136
rect 6205 1064 6211 1196
rect 6237 1064 6243 1316
rect 6253 1184 6259 1216
rect 6269 1184 6275 1196
rect 6173 1057 6195 1063
rect 6045 904 6051 996
rect 6125 944 6131 996
rect 6141 964 6147 1016
rect 6157 924 6163 1016
rect 6173 924 6179 1057
rect 6189 1024 6195 1036
rect 6189 944 6195 956
rect 5949 544 5955 556
rect 6013 504 6019 518
rect 6061 384 6067 796
rect 6109 764 6115 916
rect 6189 903 6195 916
rect 6173 897 6195 903
rect 6173 884 6179 897
rect 6205 743 6211 1016
rect 6253 1004 6259 1036
rect 6260 937 6275 943
rect 6221 784 6227 816
rect 6237 804 6243 916
rect 6269 904 6275 937
rect 6205 737 6227 743
rect 6125 684 6131 736
rect 6173 724 6179 736
rect 6141 704 6147 716
rect 6141 564 6147 576
rect 6221 524 6227 737
rect 6253 704 6259 776
rect 6269 744 6275 896
rect 6269 684 6275 736
rect 6285 724 6291 1296
rect 6317 1284 6323 1316
rect 6365 1304 6371 1336
rect 6429 1324 6435 1356
rect 6381 1144 6387 1316
rect 6429 1184 6435 1316
rect 6461 1264 6467 1356
rect 6477 1344 6483 1376
rect 6493 1324 6499 1336
rect 6461 1204 6467 1236
rect 6365 1104 6371 1116
rect 6301 924 6307 1056
rect 6333 1024 6339 1096
rect 6301 704 6307 816
rect 6317 784 6323 916
rect 6333 864 6339 936
rect 5661 224 5667 256
rect 5668 217 5683 223
rect 5677 164 5683 217
rect 5693 144 5699 236
rect 5709 204 5715 276
rect 5789 264 5795 276
rect 5821 184 5827 276
rect 5709 144 5715 156
rect 5837 144 5843 236
rect 5869 204 5875 276
rect 5885 264 5891 276
rect 5997 264 6003 316
rect 5946 214 5958 216
rect 5931 206 5933 214
rect 5941 206 5943 214
rect 5951 206 5953 214
rect 5961 206 5963 214
rect 5971 206 5973 214
rect 5946 204 5958 206
rect 5901 183 5907 196
rect 5901 177 5916 183
rect 5725 124 5731 136
rect 5997 124 6003 256
rect 6013 144 6019 336
rect 6077 284 6083 516
rect 6221 304 6227 516
rect 6253 384 6259 656
rect 6333 584 6339 856
rect 6381 703 6387 1136
rect 6461 1084 6467 1196
rect 6429 983 6435 1056
rect 6509 1024 6515 1576
rect 6589 1444 6595 1496
rect 6541 1124 6547 1436
rect 6621 1343 6627 1596
rect 6653 1564 6659 1716
rect 6669 1704 6675 1716
rect 6685 1664 6691 1736
rect 6733 1724 6739 1736
rect 6701 1584 6707 1616
rect 6765 1584 6771 1716
rect 6653 1504 6659 1556
rect 6637 1484 6643 1496
rect 6637 1384 6643 1396
rect 6653 1364 6659 1496
rect 6685 1444 6691 1496
rect 6692 1437 6707 1443
rect 6621 1337 6643 1343
rect 6589 1304 6595 1336
rect 6621 1304 6627 1316
rect 6557 1164 6563 1216
rect 6573 1184 6579 1196
rect 6541 1104 6547 1116
rect 6557 1084 6563 1156
rect 6429 977 6451 983
rect 6397 924 6403 976
rect 6429 944 6435 956
rect 6413 904 6419 916
rect 6381 697 6396 703
rect 6372 677 6396 683
rect 6365 644 6371 656
rect 6349 544 6355 576
rect 6365 344 6371 636
rect 6429 544 6435 936
rect 6445 924 6451 977
rect 6445 704 6451 856
rect 6445 584 6451 616
rect 6445 544 6451 576
rect 6461 563 6467 1016
rect 6541 937 6556 943
rect 6477 924 6483 936
rect 6493 903 6499 936
rect 6484 897 6499 903
rect 6477 724 6483 896
rect 6509 884 6515 916
rect 6525 724 6531 936
rect 6541 924 6547 937
rect 6573 924 6579 1136
rect 6637 1123 6643 1337
rect 6669 1324 6675 1396
rect 6685 1324 6691 1356
rect 6637 1117 6659 1123
rect 6605 964 6611 976
rect 6621 944 6627 956
rect 6557 903 6563 916
rect 6557 897 6579 903
rect 6573 884 6579 897
rect 6573 704 6579 856
rect 6637 763 6643 1096
rect 6621 757 6643 763
rect 6493 664 6499 696
rect 6541 644 6547 656
rect 6461 557 6483 563
rect 6381 524 6387 536
rect 6429 504 6435 516
rect 6285 304 6291 316
rect 6349 303 6355 316
rect 6333 297 6355 303
rect 6333 284 6339 297
rect 6365 284 6371 336
rect 6269 264 6275 276
rect 6093 164 6099 176
rect 6061 124 6067 136
rect 6093 124 6099 136
rect 6221 124 6227 216
rect 6397 124 6403 356
rect 6477 323 6483 557
rect 6557 544 6563 636
rect 6621 564 6627 757
rect 6541 537 6556 543
rect 6477 317 6499 323
rect 6429 302 6435 316
rect 6413 124 6419 216
rect 6477 184 6483 256
rect 6493 184 6499 317
rect 6541 244 6547 537
rect 6557 504 6563 516
rect 6653 204 6659 1117
rect 6701 1064 6707 1437
rect 6717 1324 6723 1556
rect 6765 1504 6771 1536
rect 6733 1484 6739 1496
rect 6733 1464 6739 1476
rect 6749 1444 6755 1496
rect 6781 1484 6787 2056
rect 6813 2044 6819 2116
rect 6845 2104 6851 2196
rect 6845 1904 6851 1976
rect 6861 1943 6867 2316
rect 6893 2304 6899 2676
rect 6909 2504 6915 2523
rect 6925 2284 6931 2616
rect 6941 2324 6947 3816
rect 6957 3724 6963 3836
rect 6989 3804 6995 3977
rect 7053 3884 7059 4116
rect 7085 3904 7091 4096
rect 7133 4064 7139 4276
rect 7149 3924 7155 3936
rect 7181 3924 7187 4276
rect 7197 3944 7203 4016
rect 7197 3904 7203 3936
rect 7085 3864 7091 3896
rect 7149 3884 7155 3896
rect 6973 3704 6979 3716
rect 6989 3624 6995 3636
rect 7005 3624 7011 3756
rect 7021 3664 7027 3716
rect 7021 3564 7027 3656
rect 7021 3504 7027 3516
rect 7037 3464 7043 3816
rect 7069 3784 7075 3836
rect 7053 3604 7059 3716
rect 6957 3304 6963 3316
rect 6957 3104 6963 3136
rect 6973 3084 6979 3256
rect 6989 3184 6995 3236
rect 6973 3043 6979 3076
rect 6973 3037 6995 3043
rect 6973 2944 6979 2976
rect 6989 2944 6995 3037
rect 7005 2984 7011 3456
rect 7037 3344 7043 3436
rect 7053 3324 7059 3456
rect 7037 3264 7043 3316
rect 7021 3084 7027 3116
rect 7005 2904 7011 2916
rect 6996 2877 7020 2883
rect 6973 2563 6979 2696
rect 6989 2604 6995 2676
rect 6973 2557 6995 2563
rect 6973 2484 6979 2536
rect 6925 2264 6931 2276
rect 6925 2184 6931 2196
rect 6893 2124 6899 2156
rect 6861 1937 6883 1943
rect 6845 1884 6851 1896
rect 6813 1864 6819 1876
rect 6813 1683 6819 1716
rect 6829 1704 6835 1716
rect 6813 1677 6828 1683
rect 6765 1364 6771 1396
rect 6765 1324 6771 1356
rect 6781 1324 6787 1436
rect 6797 1344 6803 1416
rect 6845 1344 6851 1536
rect 6861 1424 6867 1736
rect 6877 1544 6883 1937
rect 6893 1904 6899 2116
rect 6941 1924 6947 2176
rect 6957 1943 6963 2356
rect 6989 2164 6995 2557
rect 6957 1937 6979 1943
rect 6909 1864 6915 1896
rect 6925 1843 6931 1916
rect 6973 1884 6979 1937
rect 6909 1837 6931 1843
rect 6909 1744 6915 1837
rect 6925 1764 6931 1816
rect 6925 1704 6931 1756
rect 6925 1684 6931 1696
rect 6941 1544 6947 1636
rect 6957 1523 6963 1856
rect 6973 1744 6979 1876
rect 6989 1824 6995 1836
rect 7005 1763 7011 2596
rect 6989 1757 7011 1763
rect 6989 1724 6995 1757
rect 7021 1743 7027 2636
rect 7037 2604 7043 3096
rect 7085 3064 7091 3796
rect 7181 3764 7187 3836
rect 7117 3644 7123 3736
rect 7165 3664 7171 3696
rect 7117 3504 7123 3616
rect 7133 3524 7139 3636
rect 7181 3584 7187 3736
rect 7197 3724 7203 3736
rect 7213 3703 7219 4016
rect 7229 3944 7235 4116
rect 7277 4024 7283 4696
rect 7293 4164 7299 4276
rect 7229 3784 7235 3896
rect 7261 3884 7267 3896
rect 7229 3704 7235 3756
rect 7197 3697 7219 3703
rect 7197 3523 7203 3697
rect 7181 3517 7203 3523
rect 7117 3424 7123 3496
rect 7133 3344 7139 3376
rect 7165 3364 7171 3456
rect 7181 3384 7187 3517
rect 7213 3384 7219 3556
rect 7245 3484 7251 3636
rect 7261 3463 7267 3836
rect 7293 3784 7299 3856
rect 7357 3743 7363 4877
rect 7341 3737 7363 3743
rect 7293 3523 7299 3636
rect 7293 3517 7315 3523
rect 7245 3457 7267 3463
rect 7101 3323 7107 3336
rect 7149 3324 7155 3356
rect 7101 3317 7123 3323
rect 7117 3304 7123 3317
rect 7101 3264 7107 3296
rect 7117 2943 7123 3136
rect 7101 2937 7123 2943
rect 7085 2724 7091 2836
rect 7069 2703 7075 2716
rect 7069 2697 7084 2703
rect 7053 2124 7059 2616
rect 7101 2584 7107 2937
rect 7117 2904 7123 2916
rect 7117 2664 7123 2676
rect 7117 2564 7123 2656
rect 7133 2624 7139 3216
rect 7149 3104 7155 3176
rect 7165 2944 7171 3256
rect 7181 3084 7187 3316
rect 7197 3284 7203 3356
rect 7165 2924 7171 2936
rect 7101 2504 7107 2516
rect 7101 2224 7107 2296
rect 7117 2284 7123 2556
rect 7117 2144 7123 2276
rect 7053 1864 7059 2076
rect 7037 1764 7043 1796
rect 7012 1737 7027 1743
rect 6989 1524 6995 1536
rect 6957 1517 6979 1523
rect 6813 1324 6819 1336
rect 6717 1304 6723 1316
rect 6749 1183 6755 1276
rect 6749 1177 6764 1183
rect 6765 984 6771 1036
rect 6765 964 6771 976
rect 6749 944 6755 956
rect 6781 944 6787 1316
rect 6797 924 6803 1176
rect 6861 1104 6867 1236
rect 6829 1084 6835 1096
rect 6877 964 6883 1476
rect 6893 1404 6899 1494
rect 6957 1484 6963 1496
rect 6909 1344 6915 1416
rect 6973 1403 6979 1517
rect 6989 1504 6995 1516
rect 6957 1397 6979 1403
rect 6909 1224 6915 1336
rect 6957 1104 6963 1397
rect 6973 1104 6979 1116
rect 6957 1084 6963 1096
rect 6909 924 6915 936
rect 6708 917 6723 923
rect 6669 684 6675 876
rect 6701 783 6707 836
rect 6685 777 6707 783
rect 6685 744 6691 777
rect 6717 724 6723 917
rect 6797 864 6803 916
rect 6797 784 6803 796
rect 6813 744 6819 916
rect 6829 844 6835 916
rect 6845 784 6851 836
rect 6685 684 6691 696
rect 6749 664 6755 696
rect 6781 684 6787 696
rect 6749 544 6755 576
rect 6781 564 6787 676
rect 6797 544 6803 676
rect 6813 664 6819 736
rect 6861 704 6867 736
rect 6829 664 6835 696
rect 6877 604 6883 696
rect 6813 544 6819 556
rect 6765 504 6771 536
rect 6845 504 6851 536
rect 6781 343 6787 436
rect 6765 337 6787 343
rect 6765 324 6771 337
rect 6733 304 6739 316
rect 6829 302 6835 336
rect 6845 324 6851 496
rect 6861 284 6867 516
rect 6717 244 6723 276
rect 6861 224 6867 276
rect 6877 264 6883 596
rect 6893 544 6899 896
rect 6909 744 6915 916
rect 6925 844 6931 916
rect 6941 824 6947 836
rect 6957 764 6963 1076
rect 6973 904 6979 1096
rect 6989 944 6995 1456
rect 7005 1404 7011 1436
rect 7021 1164 7027 1576
rect 7037 1543 7043 1716
rect 7053 1684 7059 1736
rect 7053 1564 7059 1676
rect 7069 1584 7075 1896
rect 7085 1744 7091 2116
rect 7133 2103 7139 2216
rect 7149 2124 7155 2576
rect 7181 2404 7187 2436
rect 7133 2097 7155 2103
rect 7117 2084 7123 2096
rect 7101 1904 7107 1916
rect 7085 1704 7091 1716
rect 7085 1544 7091 1696
rect 7037 1537 7059 1543
rect 7053 1504 7059 1537
rect 7037 1344 7043 1496
rect 7053 1484 7059 1496
rect 7069 1424 7075 1496
rect 7085 1464 7091 1476
rect 7101 1404 7107 1856
rect 7149 1844 7155 2097
rect 7165 2084 7171 2216
rect 7181 2024 7187 2236
rect 7213 2223 7219 3356
rect 7245 3224 7251 3457
rect 7277 3324 7283 3476
rect 7309 3344 7315 3517
rect 7341 3423 7347 3737
rect 7325 3417 7347 3423
rect 7277 3163 7283 3276
rect 7293 3183 7299 3336
rect 7309 3304 7315 3316
rect 7293 3177 7315 3183
rect 7277 3157 7299 3163
rect 7245 2944 7251 3096
rect 7261 3084 7267 3156
rect 7293 3084 7299 3157
rect 7309 3104 7315 3177
rect 7309 3064 7315 3076
rect 7325 3063 7331 3417
rect 7341 3104 7347 3156
rect 7357 3064 7363 3236
rect 7325 3057 7347 3063
rect 7277 2943 7283 3036
rect 7261 2937 7283 2943
rect 7245 2684 7251 2916
rect 7245 2524 7251 2676
rect 7245 2304 7251 2516
rect 7261 2444 7267 2937
rect 7213 2217 7235 2223
rect 7181 1864 7187 1996
rect 7197 1863 7203 2176
rect 7229 2004 7235 2217
rect 7245 2124 7251 2296
rect 7245 1904 7251 2116
rect 7245 1884 7251 1896
rect 7197 1857 7219 1863
rect 7181 1824 7187 1836
rect 7133 1724 7139 1776
rect 7165 1723 7171 1756
rect 7149 1717 7171 1723
rect 7149 1624 7155 1717
rect 7181 1664 7187 1816
rect 7181 1584 7187 1616
rect 7197 1584 7203 1836
rect 7213 1803 7219 1857
rect 7213 1797 7235 1803
rect 7133 1483 7139 1496
rect 7165 1484 7171 1496
rect 7133 1477 7155 1483
rect 7133 1383 7139 1456
rect 7124 1377 7139 1383
rect 7117 1364 7123 1376
rect 7037 1304 7043 1316
rect 7053 1144 7059 1336
rect 7005 984 7011 1116
rect 7021 1044 7027 1056
rect 7028 1037 7043 1043
rect 7037 944 7043 1037
rect 7053 924 7059 976
rect 6989 784 6995 876
rect 6957 704 6963 736
rect 6925 684 6931 696
rect 6909 544 6915 576
rect 6925 564 6931 576
rect 6893 524 6899 536
rect 6957 384 6963 676
rect 6973 604 6979 696
rect 7005 463 7011 756
rect 7021 684 7027 696
rect 7053 584 7059 696
rect 7069 684 7075 696
rect 7053 524 7059 536
rect 7037 504 7043 516
rect 7005 457 7027 463
rect 7005 384 7011 436
rect 7021 284 7027 457
rect 6621 126 6627 196
rect 6157 104 6163 118
rect 6653 104 6659 136
rect 6813 126 6819 196
rect 6893 144 6899 156
rect 6845 124 6851 136
rect 6941 124 6947 156
rect 7037 144 7043 276
rect 7085 164 7091 1156
rect 7117 1104 7123 1136
rect 7101 1084 7107 1096
rect 7101 624 7107 696
rect 7117 584 7123 656
rect 7133 524 7139 1336
rect 7149 1324 7155 1477
rect 7181 1444 7187 1496
rect 7197 1143 7203 1536
rect 7213 1464 7219 1596
rect 7229 1544 7235 1797
rect 7245 1724 7251 1876
rect 7261 1683 7267 2116
rect 7277 1864 7283 2916
rect 7341 2883 7347 3057
rect 7341 2877 7363 2883
rect 7325 2684 7331 2816
rect 7357 2704 7363 2877
rect 7373 2703 7379 3516
rect 7405 3324 7411 4536
rect 7389 3024 7395 3056
rect 7373 2697 7395 2703
rect 7341 2184 7347 2636
rect 7373 2584 7379 2676
rect 7277 1764 7283 1836
rect 7277 1704 7283 1716
rect 7261 1677 7283 1683
rect 7277 1584 7283 1677
rect 7181 1137 7203 1143
rect 7149 944 7155 1056
rect 7165 924 7171 976
rect 7149 604 7155 656
rect 7181 603 7187 1137
rect 7213 1084 7219 1336
rect 7245 1104 7251 1116
rect 7213 924 7219 1056
rect 7229 984 7235 1076
rect 7245 964 7251 1096
rect 7245 944 7251 956
rect 7261 924 7267 1056
rect 7229 784 7235 876
rect 7229 704 7235 736
rect 7165 597 7187 603
rect 7149 544 7155 556
rect 7165 504 7171 597
rect 7245 564 7251 896
rect 7277 884 7283 1556
rect 7293 1504 7299 2096
rect 7341 1784 7347 2016
rect 7293 1484 7299 1496
rect 7325 1464 7331 1776
rect 7357 1584 7363 1836
rect 7341 1344 7347 1396
rect 7309 1304 7315 1336
rect 7293 1084 7299 1116
rect 7293 983 7299 1016
rect 7309 1004 7315 1096
rect 7325 1084 7331 1236
rect 7357 1084 7363 1536
rect 7373 1484 7379 1816
rect 7357 1064 7363 1076
rect 7325 984 7331 1056
rect 7341 984 7347 1036
rect 7293 977 7315 983
rect 7261 724 7267 816
rect 7293 804 7299 956
rect 7309 944 7315 977
rect 7341 944 7347 956
rect 7309 704 7315 916
rect 7245 284 7251 516
rect 7261 364 7267 696
rect 7309 684 7315 696
rect 7325 644 7331 696
rect 7341 683 7347 936
rect 7357 824 7363 1036
rect 7357 784 7363 796
rect 7373 704 7379 956
rect 7341 677 7363 683
rect 7293 524 7299 616
rect 7357 583 7363 677
rect 7341 577 7363 583
rect 7341 383 7347 577
rect 7341 377 7356 383
rect 7389 204 7395 2697
rect 7405 1804 7411 2756
rect 7069 104 7075 116
rect 5149 97 5164 103
rect 5149 -23 5155 97
rect 5213 23 5219 96
rect 5204 17 5219 23
rect 5197 -23 5203 16
<< m3contact >>
rect 1036 5396 1044 5404
rect 1100 5396 1108 5404
rect 460 5376 468 5384
rect 508 5376 516 5384
rect 316 5356 324 5364
rect 396 5356 404 5364
rect 44 5316 52 5324
rect 156 5316 164 5324
rect 204 5316 212 5324
rect 12 5296 20 5304
rect 108 5296 116 5304
rect 284 5336 292 5344
rect 364 5336 372 5344
rect 380 5336 388 5344
rect 428 5336 436 5344
rect 620 5356 628 5364
rect 796 5356 804 5364
rect 844 5356 852 5364
rect 956 5356 964 5364
rect 492 5336 500 5344
rect 540 5336 548 5344
rect 572 5336 580 5344
rect 748 5336 756 5344
rect 764 5336 772 5344
rect 796 5336 804 5344
rect 252 5256 260 5264
rect 140 5136 148 5144
rect 12 5096 20 5104
rect 60 5096 68 5104
rect 108 5096 116 5104
rect 156 5096 164 5104
rect 188 5096 196 5104
rect 236 5096 244 5104
rect 236 5076 244 5084
rect 316 5216 324 5224
rect 300 5096 308 5104
rect 76 5056 84 5064
rect 124 5056 132 5064
rect 220 5056 228 5064
rect 252 5056 260 5064
rect 300 5056 308 5064
rect 76 5036 84 5044
rect 60 4976 68 4984
rect 140 4936 148 4944
rect 12 4736 20 4744
rect 44 4736 52 4744
rect 204 4976 212 4984
rect 252 4976 260 4984
rect 204 4956 212 4964
rect 332 5096 340 5104
rect 524 5116 532 5124
rect 380 5096 388 5104
rect 412 5096 420 5104
rect 396 5076 404 5084
rect 444 5076 452 5084
rect 652 5316 660 5324
rect 652 5276 660 5284
rect 700 5316 708 5324
rect 764 5316 772 5324
rect 668 5256 676 5264
rect 748 5256 756 5264
rect 908 5316 916 5324
rect 1004 5316 1012 5324
rect 844 5256 852 5264
rect 892 5256 900 5264
rect 972 5256 980 5264
rect 812 5236 820 5244
rect 556 5116 564 5124
rect 604 5116 612 5124
rect 636 5116 644 5124
rect 684 5116 692 5124
rect 556 5096 564 5104
rect 588 5096 596 5104
rect 540 5076 548 5084
rect 428 5056 436 5064
rect 492 5056 500 5064
rect 348 5036 356 5044
rect 252 4936 260 4944
rect 172 4916 180 4924
rect 220 4916 228 4924
rect 124 4736 132 4744
rect 140 4736 148 4744
rect 204 4736 212 4744
rect 156 4716 164 4724
rect 156 4676 164 4684
rect 76 4556 84 4564
rect 124 4556 132 4564
rect 236 4756 244 4764
rect 492 5016 500 5024
rect 396 4976 404 4984
rect 524 4996 532 5004
rect 492 4936 500 4944
rect 508 4936 516 4944
rect 364 4916 372 4924
rect 412 4916 420 4924
rect 636 5096 644 5104
rect 748 5096 756 5104
rect 796 5096 804 5104
rect 668 5056 676 5064
rect 604 4996 612 5004
rect 860 5176 868 5184
rect 972 5136 980 5144
rect 828 5096 836 5104
rect 716 5076 724 5084
rect 812 5076 820 5084
rect 732 5056 740 5064
rect 828 5056 836 5064
rect 956 5096 964 5104
rect 892 5056 900 5064
rect 860 5036 868 5044
rect 684 4976 692 4984
rect 540 4956 548 4964
rect 588 4956 596 4964
rect 604 4956 612 4964
rect 684 4956 692 4964
rect 716 4956 724 4964
rect 588 4936 596 4944
rect 620 4936 628 4944
rect 668 4936 676 4944
rect 316 4896 324 4904
rect 284 4696 292 4704
rect 332 4696 340 4704
rect 236 4656 244 4664
rect 284 4656 292 4664
rect 220 4616 228 4624
rect 572 4916 580 4924
rect 732 4916 740 4924
rect 476 4876 484 4884
rect 636 4876 644 4884
rect 764 4896 772 4904
rect 428 4796 436 4804
rect 508 4756 516 4764
rect 556 4756 564 4764
rect 588 4756 596 4764
rect 364 4736 372 4744
rect 460 4716 468 4724
rect 428 4696 436 4704
rect 460 4656 468 4664
rect 348 4636 356 4644
rect 396 4616 404 4624
rect 268 4576 276 4584
rect 316 4576 324 4584
rect 332 4576 340 4584
rect 140 4536 148 4544
rect 188 4536 196 4544
rect 572 4696 580 4704
rect 732 4736 740 4744
rect 620 4696 628 4704
rect 796 4716 804 4724
rect 908 4956 916 4964
rect 892 4716 900 4724
rect 844 4696 852 4704
rect 812 4676 820 4684
rect 636 4656 644 4664
rect 668 4656 676 4664
rect 508 4636 516 4644
rect 492 4616 500 4624
rect 444 4576 452 4584
rect 476 4576 484 4584
rect 428 4556 436 4564
rect 492 4556 500 4564
rect 396 4536 404 4544
rect 476 4536 484 4544
rect 12 4516 20 4524
rect 44 4516 52 4524
rect 92 4516 100 4524
rect 204 4516 212 4524
rect 300 4516 308 4524
rect 28 4496 36 4504
rect 92 4496 100 4504
rect 124 4336 132 4344
rect 108 4276 116 4284
rect 140 4316 148 4324
rect 460 4496 468 4504
rect 364 4476 372 4484
rect 236 4336 244 4344
rect 268 4336 276 4344
rect 172 4276 180 4284
rect 284 4296 292 4304
rect 44 4256 52 4264
rect 140 4256 148 4264
rect 220 4256 228 4264
rect 60 4196 68 4204
rect 236 4196 244 4204
rect 44 4116 52 4124
rect 108 4176 116 4184
rect 156 4156 164 4164
rect 76 4116 84 4124
rect 140 4096 148 4104
rect 28 4076 36 4084
rect 92 4076 100 4084
rect 12 3956 20 3964
rect 12 3936 20 3944
rect 44 3936 52 3944
rect 44 3916 52 3924
rect 124 3916 132 3924
rect 316 4256 324 4264
rect 220 4096 228 4104
rect 204 4036 212 4044
rect 236 4036 244 4044
rect 252 3916 260 3924
rect 60 3896 68 3904
rect 124 3896 132 3904
rect 156 3896 164 3904
rect 236 3896 244 3904
rect 12 3756 20 3764
rect 28 3476 36 3484
rect 108 3876 116 3884
rect 236 3876 244 3884
rect 188 3836 196 3844
rect 220 3836 228 3844
rect 188 3816 196 3824
rect 284 3876 292 3884
rect 268 3856 276 3864
rect 300 3856 308 3864
rect 636 4596 644 4604
rect 524 4556 532 4564
rect 588 4556 596 4564
rect 524 4496 532 4504
rect 572 4476 580 4484
rect 508 4396 516 4404
rect 348 4336 356 4344
rect 364 4316 372 4324
rect 396 4296 404 4304
rect 604 4356 612 4364
rect 716 4616 724 4624
rect 700 4596 708 4604
rect 716 4576 724 4584
rect 684 4536 692 4544
rect 764 4596 772 4604
rect 812 4656 820 4664
rect 812 4616 820 4624
rect 844 4576 852 4584
rect 828 4556 836 4564
rect 764 4536 772 4544
rect 844 4516 852 4524
rect 652 4376 660 4384
rect 620 4336 628 4344
rect 668 4336 676 4344
rect 556 4316 564 4324
rect 620 4316 628 4324
rect 748 4316 756 4324
rect 876 4696 884 4704
rect 2556 5416 2564 5424
rect 1324 5376 1332 5384
rect 1484 5376 1492 5384
rect 1916 5376 1924 5384
rect 2028 5376 2036 5384
rect 2284 5376 2292 5384
rect 2332 5376 2340 5384
rect 1084 5356 1092 5364
rect 1212 5356 1220 5364
rect 1276 5356 1284 5364
rect 1564 5356 1572 5364
rect 1644 5356 1652 5364
rect 1836 5356 1844 5364
rect 1900 5356 1908 5364
rect 1068 5336 1076 5344
rect 1052 5316 1060 5324
rect 1180 5316 1188 5324
rect 1132 5256 1140 5264
rect 1020 5236 1028 5244
rect 1180 5296 1188 5304
rect 1164 5216 1172 5224
rect 1116 5176 1124 5184
rect 1100 5156 1108 5164
rect 1036 5096 1044 5104
rect 1052 5096 1060 5104
rect 1100 5096 1108 5104
rect 1004 5076 1012 5084
rect 1148 5156 1156 5164
rect 1164 5156 1172 5164
rect 1356 5256 1364 5264
rect 1324 5176 1332 5184
rect 1164 5136 1172 5144
rect 1228 5136 1236 5144
rect 1148 5096 1156 5104
rect 1164 5096 1172 5104
rect 1196 5096 1204 5104
rect 1212 5096 1220 5104
rect 1260 5096 1268 5104
rect 1308 5096 1316 5104
rect 1036 5076 1044 5084
rect 1132 5076 1140 5084
rect 1596 5336 1604 5344
rect 1500 5296 1508 5304
rect 1372 5236 1380 5244
rect 1404 5236 1412 5244
rect 1411 5206 1419 5214
rect 1421 5206 1429 5214
rect 1431 5206 1439 5214
rect 1441 5206 1449 5214
rect 1451 5206 1459 5214
rect 1461 5206 1469 5214
rect 1436 5136 1444 5144
rect 1484 5136 1492 5144
rect 1212 5076 1220 5084
rect 1020 5056 1028 5064
rect 1004 5016 1012 5024
rect 988 4956 996 4964
rect 940 4936 948 4944
rect 988 4936 996 4944
rect 1068 5016 1076 5024
rect 1292 5056 1300 5064
rect 1340 5056 1348 5064
rect 1244 4996 1252 5004
rect 1356 4996 1364 5004
rect 1292 4976 1300 4984
rect 1308 4976 1316 4984
rect 1148 4956 1156 4964
rect 1068 4936 1076 4944
rect 940 4916 948 4924
rect 972 4916 980 4924
rect 1004 4916 1012 4924
rect 1036 4916 1044 4924
rect 924 4896 932 4904
rect 1164 4936 1172 4944
rect 1196 4936 1204 4944
rect 1228 4956 1236 4964
rect 1260 4956 1268 4964
rect 1116 4916 1124 4924
rect 1244 4916 1252 4924
rect 1276 4936 1284 4944
rect 1324 4916 1332 4924
rect 1260 4876 1268 4884
rect 1324 4876 1332 4884
rect 1340 4876 1348 4884
rect 1100 4776 1108 4784
rect 1052 4756 1060 4764
rect 1100 4756 1108 4764
rect 988 4736 996 4744
rect 1052 4736 1060 4744
rect 1004 4716 1012 4724
rect 1084 4716 1092 4724
rect 956 4676 964 4684
rect 908 4656 916 4664
rect 940 4636 948 4644
rect 1004 4636 1012 4644
rect 1068 4636 1076 4644
rect 892 4556 900 4564
rect 924 4556 932 4564
rect 1052 4616 1060 4624
rect 1116 4736 1124 4744
rect 1100 4676 1108 4684
rect 1180 4676 1188 4684
rect 1116 4656 1124 4664
rect 1020 4576 1028 4584
rect 1084 4576 1092 4584
rect 892 4516 900 4524
rect 1164 4596 1172 4604
rect 1132 4556 1140 4564
rect 1372 4936 1380 4944
rect 1372 4876 1380 4884
rect 1596 5296 1604 5304
rect 1628 5336 1636 5344
rect 1692 5336 1700 5344
rect 1660 5296 1668 5304
rect 1612 5256 1620 5264
rect 1596 5136 1604 5144
rect 1516 5096 1524 5104
rect 1548 5096 1556 5104
rect 1692 5256 1700 5264
rect 1964 5356 1972 5364
rect 1996 5356 2004 5364
rect 1852 5316 1860 5324
rect 1916 5316 1924 5324
rect 1932 5316 1940 5324
rect 1788 5296 1796 5304
rect 1804 5296 1812 5304
rect 1708 5236 1716 5244
rect 1756 5236 1764 5244
rect 1820 5196 1828 5204
rect 1804 5176 1812 5184
rect 1820 5176 1828 5184
rect 1660 5096 1668 5104
rect 1772 5096 1780 5104
rect 1788 5096 1796 5104
rect 1932 5296 1940 5304
rect 1980 5296 1988 5304
rect 1916 5176 1924 5184
rect 1868 5156 1876 5164
rect 1836 5136 1844 5144
rect 1516 4976 1524 4984
rect 1420 4956 1428 4964
rect 1436 4956 1444 4964
rect 1500 4956 1508 4964
rect 1532 4956 1540 4964
rect 1516 4936 1524 4944
rect 1580 4936 1588 4944
rect 1644 5036 1652 5044
rect 1692 5076 1700 5084
rect 1708 5076 1716 5084
rect 1724 5076 1732 5084
rect 1804 5076 1812 5084
rect 1676 5056 1684 5064
rect 1692 5056 1700 5064
rect 1612 4956 1620 4964
rect 1404 4856 1412 4864
rect 1420 4856 1428 4864
rect 1532 4836 1540 4844
rect 1411 4806 1419 4814
rect 1421 4806 1429 4814
rect 1431 4806 1439 4814
rect 1441 4806 1449 4814
rect 1451 4806 1459 4814
rect 1461 4806 1469 4814
rect 1468 4776 1476 4784
rect 1356 4736 1364 4744
rect 1308 4716 1316 4724
rect 1356 4716 1364 4724
rect 1260 4696 1268 4704
rect 1276 4696 1284 4704
rect 1372 4696 1380 4704
rect 1292 4676 1300 4684
rect 1340 4656 1348 4664
rect 1212 4596 1220 4604
rect 1196 4576 1204 4584
rect 1308 4616 1316 4624
rect 1052 4516 1060 4524
rect 1084 4516 1092 4524
rect 956 4496 964 4504
rect 1132 4496 1140 4504
rect 700 4296 708 4304
rect 492 4276 500 4284
rect 604 4276 612 4284
rect 652 4276 660 4284
rect 380 4256 388 4264
rect 364 4236 372 4244
rect 428 4256 436 4264
rect 508 4256 516 4264
rect 604 4256 612 4264
rect 412 4236 420 4244
rect 620 4236 628 4244
rect 668 4236 676 4244
rect 460 4196 468 4204
rect 460 4176 468 4184
rect 924 4376 932 4384
rect 988 4336 996 4344
rect 892 4316 900 4324
rect 972 4316 980 4324
rect 748 4276 756 4284
rect 1148 4396 1156 4404
rect 1148 4336 1156 4344
rect 1068 4316 1076 4324
rect 1052 4296 1060 4304
rect 924 4276 932 4284
rect 860 4236 868 4244
rect 892 4236 900 4244
rect 780 4216 788 4224
rect 700 4196 708 4204
rect 700 4176 708 4184
rect 540 4156 548 4164
rect 524 4136 532 4144
rect 428 4016 436 4024
rect 396 3936 404 3944
rect 348 3916 356 3924
rect 540 3916 548 3924
rect 460 3896 468 3904
rect 476 3896 484 3904
rect 364 3876 372 3884
rect 460 3856 468 3864
rect 332 3836 340 3844
rect 316 3816 324 3824
rect 60 3756 68 3764
rect 252 3756 260 3764
rect 524 3876 532 3884
rect 428 3776 436 3784
rect 476 3776 484 3784
rect 540 3856 548 3864
rect 604 4036 612 4044
rect 732 4136 740 4144
rect 828 4156 836 4164
rect 812 4136 820 4144
rect 844 4116 852 4124
rect 636 4016 644 4024
rect 620 3936 628 3944
rect 684 3936 692 3944
rect 572 3916 580 3924
rect 652 3916 660 3924
rect 700 3916 708 3924
rect 716 3876 724 3884
rect 572 3856 580 3864
rect 652 3856 660 3864
rect 716 3856 724 3864
rect 732 3816 740 3824
rect 460 3756 468 3764
rect 524 3756 532 3764
rect 556 3756 564 3764
rect 716 3756 724 3764
rect 236 3736 244 3744
rect 284 3736 292 3744
rect 396 3736 404 3744
rect 412 3736 420 3744
rect 476 3736 484 3744
rect 556 3736 564 3744
rect 108 3716 116 3724
rect 156 3716 164 3724
rect 508 3716 516 3724
rect 604 3716 612 3724
rect 668 3716 676 3724
rect 60 3576 68 3584
rect 92 3496 100 3504
rect 108 3476 116 3484
rect 44 3336 52 3344
rect 124 3336 132 3344
rect 140 3316 148 3324
rect 108 3296 116 3304
rect 140 3296 148 3304
rect 396 3696 404 3704
rect 428 3696 436 3704
rect 316 3676 324 3684
rect 172 3576 180 3584
rect 284 3576 292 3584
rect 332 3536 340 3544
rect 220 3496 228 3504
rect 252 3496 260 3504
rect 316 3496 324 3504
rect 172 3456 180 3464
rect 204 3456 212 3464
rect 172 3416 180 3424
rect 172 3276 180 3284
rect 108 3136 116 3144
rect 92 3076 100 3084
rect 76 3056 84 3064
rect 92 2916 100 2924
rect 156 2916 164 2924
rect 92 2696 100 2704
rect 60 2516 68 2524
rect 300 3476 308 3484
rect 284 3356 292 3364
rect 588 3696 596 3704
rect 588 3636 596 3644
rect 620 3636 628 3644
rect 556 3576 564 3584
rect 412 3536 420 3544
rect 460 3536 468 3544
rect 508 3536 516 3544
rect 428 3476 436 3484
rect 572 3476 580 3484
rect 684 3596 692 3604
rect 700 3496 708 3504
rect 732 3596 740 3604
rect 780 3916 788 3924
rect 764 3896 772 3904
rect 764 3816 772 3824
rect 988 4196 996 4204
rect 1052 4216 1060 4224
rect 1004 4176 1012 4184
rect 1020 4176 1028 4184
rect 1036 4176 1044 4184
rect 1052 4176 1060 4184
rect 924 4156 932 4164
rect 940 4156 948 4164
rect 1132 4236 1140 4244
rect 1116 4196 1124 4204
rect 956 4136 964 4144
rect 1084 4136 1092 4144
rect 972 4116 980 4124
rect 1020 4116 1028 4124
rect 1084 4116 1092 4124
rect 1052 4096 1060 4104
rect 1004 4076 1012 4084
rect 1132 4076 1140 4084
rect 908 4056 916 4064
rect 876 4036 884 4044
rect 860 3996 868 4004
rect 860 3936 868 3944
rect 812 3916 820 3924
rect 908 4016 916 4024
rect 892 3956 900 3964
rect 844 3876 852 3884
rect 876 3856 884 3864
rect 812 3816 820 3824
rect 828 3816 836 3824
rect 780 3756 788 3764
rect 860 3836 868 3844
rect 844 3756 852 3764
rect 1036 3916 1044 3924
rect 924 3896 932 3904
rect 1100 3996 1108 4004
rect 1132 4036 1140 4044
rect 908 3796 916 3804
rect 844 3716 852 3724
rect 908 3716 916 3724
rect 828 3676 836 3684
rect 812 3616 820 3624
rect 748 3556 756 3564
rect 796 3556 804 3564
rect 812 3496 820 3504
rect 556 3456 564 3464
rect 268 3336 276 3344
rect 332 3336 340 3344
rect 492 3396 500 3404
rect 492 3376 500 3384
rect 428 3336 436 3344
rect 460 3296 468 3304
rect 524 3356 532 3364
rect 556 3356 564 3364
rect 508 3296 516 3304
rect 412 3156 420 3164
rect 348 3136 356 3144
rect 252 3116 260 3124
rect 332 3116 340 3124
rect 204 3096 212 3104
rect 268 3076 276 3084
rect 252 3056 260 3064
rect 300 3056 308 3064
rect 204 3036 212 3044
rect 188 2956 196 2964
rect 268 2956 276 2964
rect 284 2936 292 2944
rect 204 2916 212 2924
rect 236 2856 244 2864
rect 204 2836 212 2844
rect 284 2856 292 2864
rect 252 2836 260 2844
rect 236 2656 244 2664
rect 108 2496 116 2504
rect 108 2316 116 2324
rect 140 2296 148 2304
rect 92 2276 100 2284
rect 12 2256 20 2264
rect 124 2256 132 2264
rect 44 2116 52 2124
rect 92 2076 100 2084
rect 140 2056 148 2064
rect 60 1916 68 1924
rect 108 1896 116 1904
rect 12 1876 20 1884
rect 108 1876 116 1884
rect 140 1876 148 1884
rect 140 1856 148 1864
rect 204 2536 212 2544
rect 236 2536 244 2544
rect 204 2516 212 2524
rect 204 2136 212 2144
rect 172 2096 180 2104
rect 172 2076 180 2084
rect 252 2496 260 2504
rect 236 2316 244 2324
rect 300 2696 308 2704
rect 364 3096 372 3104
rect 364 3056 372 3064
rect 364 2936 372 2944
rect 380 2876 388 2884
rect 412 3056 420 3064
rect 476 3056 484 3064
rect 508 3056 516 3064
rect 460 3036 468 3044
rect 412 2936 420 2944
rect 492 2956 500 2964
rect 396 2836 404 2844
rect 348 2816 356 2824
rect 332 2676 340 2684
rect 332 2656 340 2664
rect 316 2636 324 2644
rect 396 2736 404 2744
rect 428 2876 436 2884
rect 476 2916 484 2924
rect 492 2816 500 2824
rect 460 2756 468 2764
rect 444 2736 452 2744
rect 364 2616 372 2624
rect 396 2556 404 2564
rect 316 2536 324 2544
rect 380 2536 388 2544
rect 460 2536 468 2544
rect 332 2476 340 2484
rect 396 2476 404 2484
rect 444 2476 452 2484
rect 284 2296 292 2304
rect 268 2156 276 2164
rect 380 2336 388 2344
rect 428 2336 436 2344
rect 524 2816 532 2824
rect 508 2776 516 2784
rect 508 2716 516 2724
rect 508 2536 516 2544
rect 556 3096 564 3104
rect 588 3076 596 3084
rect 556 3056 564 3064
rect 620 3356 628 3364
rect 620 3316 628 3324
rect 652 3396 660 3404
rect 636 3296 644 3304
rect 620 3096 628 3104
rect 764 3476 772 3484
rect 748 3456 756 3464
rect 780 3396 788 3404
rect 812 3396 820 3404
rect 796 3356 804 3364
rect 668 3316 676 3324
rect 700 3316 708 3324
rect 764 3316 772 3324
rect 812 3316 820 3324
rect 668 3276 676 3284
rect 732 3276 740 3284
rect 700 3216 708 3224
rect 684 3116 692 3124
rect 764 3256 772 3264
rect 748 3236 756 3244
rect 764 3196 772 3204
rect 748 3116 756 3124
rect 668 3076 676 3084
rect 732 3076 740 3084
rect 812 3156 820 3164
rect 796 3136 804 3144
rect 780 3076 788 3084
rect 732 3056 740 3064
rect 764 3056 772 3064
rect 636 3036 644 3044
rect 604 2956 612 2964
rect 620 2956 628 2964
rect 572 2936 580 2944
rect 604 2916 612 2924
rect 572 2876 580 2884
rect 636 2916 644 2924
rect 716 2956 724 2964
rect 764 2976 772 2984
rect 684 2916 692 2924
rect 748 2916 756 2924
rect 668 2876 676 2884
rect 668 2836 676 2844
rect 652 2756 660 2764
rect 588 2736 596 2744
rect 620 2736 628 2744
rect 764 2876 772 2884
rect 716 2856 724 2864
rect 700 2796 708 2804
rect 780 2796 788 2804
rect 812 3096 820 3104
rect 812 2916 820 2924
rect 876 3696 884 3704
rect 1020 3856 1028 3864
rect 1068 3856 1076 3864
rect 972 3816 980 3824
rect 940 3756 948 3764
rect 988 3776 996 3784
rect 1036 3776 1044 3784
rect 1116 3896 1124 3904
rect 1148 4016 1156 4024
rect 1180 4496 1188 4504
rect 1228 4316 1236 4324
rect 1180 4296 1188 4304
rect 1228 4296 1236 4304
rect 1260 4296 1268 4304
rect 1212 4276 1220 4284
rect 1180 4256 1188 4264
rect 1196 4236 1204 4244
rect 1180 4136 1188 4144
rect 1164 3996 1172 4004
rect 1180 3936 1188 3944
rect 1228 4216 1236 4224
rect 1324 4536 1332 4544
rect 1324 4356 1332 4364
rect 1292 4316 1300 4324
rect 1596 4916 1604 4924
rect 1772 5016 1780 5024
rect 1756 4996 1764 5004
rect 1836 5096 1844 5104
rect 1852 5076 1860 5084
rect 1820 4976 1828 4984
rect 1804 4956 1812 4964
rect 1868 5016 1876 5024
rect 1852 4956 1860 4964
rect 1932 5136 1940 5144
rect 1900 5056 1908 5064
rect 1900 4956 1908 4964
rect 1836 4936 1844 4944
rect 1868 4936 1876 4944
rect 1756 4916 1764 4924
rect 2076 5356 2084 5364
rect 2108 5356 2116 5364
rect 2204 5356 2212 5364
rect 2380 5356 2388 5364
rect 2524 5336 2532 5344
rect 2044 5316 2052 5324
rect 2204 5316 2212 5324
rect 2092 5296 2100 5304
rect 2092 5256 2100 5264
rect 2012 5236 2020 5244
rect 2012 5176 2020 5184
rect 2044 5176 2052 5184
rect 2108 5196 2116 5204
rect 2268 5316 2276 5324
rect 2316 5316 2324 5324
rect 2364 5316 2372 5324
rect 2428 5316 2436 5324
rect 2220 5296 2228 5304
rect 2172 5276 2180 5284
rect 2156 5256 2164 5264
rect 2524 5296 2532 5304
rect 2268 5196 2276 5204
rect 2268 5176 2276 5184
rect 2364 5176 2372 5184
rect 2108 5076 2116 5084
rect 2156 5076 2164 5084
rect 2108 5056 2116 5064
rect 1996 5016 2004 5024
rect 1964 4956 1972 4964
rect 1996 4936 2004 4944
rect 1964 4916 1972 4924
rect 1980 4916 1988 4924
rect 2044 5016 2052 5024
rect 2076 4976 2084 4984
rect 2076 4956 2084 4964
rect 1980 4856 1988 4864
rect 2028 4856 2036 4864
rect 1660 4836 1668 4844
rect 1836 4836 1844 4844
rect 1868 4836 1876 4844
rect 1612 4816 1620 4824
rect 1580 4736 1588 4744
rect 1932 4816 1940 4824
rect 1612 4696 1620 4704
rect 1724 4696 1732 4704
rect 1788 4696 1796 4704
rect 1836 4696 1844 4704
rect 1516 4676 1524 4684
rect 1388 4656 1396 4664
rect 1580 4656 1588 4664
rect 1372 4540 1380 4544
rect 1372 4536 1380 4540
rect 1404 4536 1412 4544
rect 1372 4476 1380 4484
rect 1356 4336 1364 4344
rect 1468 4516 1476 4524
rect 1411 4406 1419 4414
rect 1421 4406 1429 4414
rect 1431 4406 1439 4414
rect 1441 4406 1449 4414
rect 1451 4406 1459 4414
rect 1461 4406 1469 4414
rect 1388 4376 1396 4384
rect 1420 4376 1428 4384
rect 1436 4356 1444 4364
rect 1516 4516 1524 4524
rect 1596 4636 1604 4644
rect 1564 4596 1572 4604
rect 1660 4636 1668 4644
rect 1724 4636 1732 4644
rect 1564 4536 1572 4544
rect 1612 4536 1620 4544
rect 1628 4536 1636 4544
rect 1756 4676 1764 4684
rect 1772 4656 1780 4664
rect 1804 4656 1812 4664
rect 1932 4656 1940 4664
rect 1852 4636 1860 4644
rect 1756 4596 1764 4604
rect 1916 4596 1924 4604
rect 1708 4556 1716 4564
rect 1740 4556 1748 4564
rect 1964 4676 1972 4684
rect 1948 4616 1956 4624
rect 2012 4736 2020 4744
rect 1996 4696 2004 4704
rect 1996 4656 2004 4664
rect 1980 4576 1988 4584
rect 1548 4496 1556 4504
rect 1500 4376 1508 4384
rect 1372 4296 1380 4304
rect 1484 4336 1492 4344
rect 1324 4276 1332 4284
rect 1372 4276 1380 4284
rect 1308 4256 1316 4264
rect 1276 4216 1284 4224
rect 1308 4156 1316 4164
rect 1276 4116 1284 4124
rect 1340 4116 1348 4124
rect 1404 4216 1412 4224
rect 1436 4196 1444 4204
rect 1436 4136 1444 4144
rect 1276 4056 1284 4064
rect 1692 4496 1700 4504
rect 1772 4476 1780 4484
rect 1612 4376 1620 4384
rect 1660 4356 1668 4364
rect 1628 4336 1636 4344
rect 1532 4296 1540 4304
rect 1692 4336 1700 4344
rect 1740 4296 1748 4304
rect 1724 4276 1732 4284
rect 1740 4256 1748 4264
rect 1708 4236 1716 4244
rect 1756 4236 1764 4244
rect 1644 4216 1652 4224
rect 1708 4156 1716 4164
rect 1788 4336 1796 4344
rect 2028 4696 2036 4704
rect 2172 4996 2180 5004
rect 2204 5136 2212 5144
rect 2476 5136 2484 5144
rect 2284 5116 2292 5124
rect 2348 5116 2356 5124
rect 2428 5116 2436 5124
rect 2460 5116 2468 5124
rect 2236 5096 2244 5104
rect 2220 4996 2228 5004
rect 2300 5076 2308 5084
rect 2380 5076 2388 5084
rect 2444 5076 2452 5084
rect 2268 5036 2276 5044
rect 2156 4936 2164 4944
rect 2252 4956 2260 4964
rect 2332 4996 2340 5004
rect 2300 4956 2308 4964
rect 2364 4956 2372 4964
rect 2460 4956 2468 4964
rect 2588 5416 2596 5424
rect 2915 5406 2923 5414
rect 2925 5406 2933 5414
rect 2935 5406 2943 5414
rect 2945 5406 2953 5414
rect 2955 5406 2963 5414
rect 2965 5406 2973 5414
rect 2684 5356 2692 5364
rect 2588 5336 2596 5344
rect 2748 5336 2756 5344
rect 2716 5318 2724 5324
rect 2716 5316 2724 5318
rect 2556 5296 2564 5304
rect 2684 5296 2692 5304
rect 2604 5076 2612 5084
rect 2540 5056 2548 5064
rect 2588 5016 2596 5024
rect 2540 4996 2548 5004
rect 2492 4976 2500 4984
rect 2636 4996 2644 5004
rect 2620 4976 2628 4984
rect 2380 4936 2388 4944
rect 2476 4936 2484 4944
rect 2508 4936 2516 4944
rect 2524 4936 2532 4944
rect 2588 4936 2596 4944
rect 2092 4916 2100 4924
rect 2124 4916 2132 4924
rect 2156 4916 2164 4924
rect 2236 4916 2244 4924
rect 2412 4916 2420 4924
rect 2476 4916 2484 4924
rect 2428 4876 2436 4884
rect 2316 4856 2324 4864
rect 2556 4856 2564 4864
rect 2332 4836 2340 4844
rect 2460 4836 2468 4844
rect 2508 4836 2516 4844
rect 2076 4816 2084 4824
rect 2204 4796 2212 4804
rect 2300 4776 2308 4784
rect 2060 4736 2068 4744
rect 2140 4736 2148 4744
rect 2204 4736 2212 4744
rect 2108 4716 2116 4724
rect 2092 4696 2100 4704
rect 2060 4636 2068 4644
rect 2076 4636 2084 4644
rect 2220 4696 2228 4704
rect 2300 4696 2308 4704
rect 2316 4696 2324 4704
rect 2172 4676 2180 4684
rect 2156 4656 2164 4664
rect 2204 4636 2212 4644
rect 2156 4576 2164 4584
rect 2220 4576 2228 4584
rect 2236 4576 2244 4584
rect 2076 4556 2084 4564
rect 2140 4556 2148 4564
rect 2012 4536 2020 4544
rect 2124 4536 2132 4544
rect 1900 4496 1908 4504
rect 2204 4556 2212 4564
rect 1932 4496 1940 4504
rect 1948 4476 1956 4484
rect 1916 4436 1924 4444
rect 1868 4356 1876 4364
rect 1900 4336 1908 4344
rect 1932 4296 1940 4304
rect 1820 4276 1828 4284
rect 1884 4276 1892 4284
rect 1916 4276 1924 4284
rect 1820 4256 1828 4264
rect 1868 4256 1876 4264
rect 1836 4236 1844 4244
rect 1596 4136 1604 4144
rect 1484 4016 1492 4024
rect 1411 4006 1419 4014
rect 1421 4006 1429 4014
rect 1431 4006 1439 4014
rect 1441 4006 1449 4014
rect 1451 4006 1459 4014
rect 1461 4006 1469 4014
rect 1388 3996 1396 4004
rect 1372 3936 1380 3944
rect 1820 4156 1828 4164
rect 1580 4116 1588 4124
rect 1692 4116 1700 4124
rect 1660 4096 1668 4104
rect 1740 4096 1748 4104
rect 1852 4096 1860 4104
rect 1580 4076 1588 4084
rect 1468 3936 1476 3944
rect 1532 3936 1540 3944
rect 1196 3896 1204 3904
rect 1260 3896 1268 3904
rect 1276 3896 1284 3904
rect 1388 3896 1396 3904
rect 1260 3836 1268 3844
rect 1324 3836 1332 3844
rect 1100 3776 1108 3784
rect 1180 3736 1188 3744
rect 1244 3736 1252 3744
rect 1564 3896 1572 3904
rect 1964 4416 1972 4424
rect 1996 4516 2004 4524
rect 2060 4516 2068 4524
rect 2044 4496 2052 4504
rect 1996 4456 2004 4464
rect 1980 4376 1988 4384
rect 1980 4356 1988 4364
rect 1964 4196 1972 4204
rect 1948 4176 1956 4184
rect 1900 4136 1908 4144
rect 1980 4156 1988 4164
rect 2028 4436 2036 4444
rect 2428 4796 2436 4804
rect 2364 4716 2372 4724
rect 2396 4696 2404 4704
rect 2492 4796 2500 4804
rect 2508 4796 2516 4804
rect 2412 4676 2420 4684
rect 2540 4736 2548 4744
rect 2380 4656 2388 4664
rect 2364 4636 2372 4644
rect 2316 4576 2324 4584
rect 2316 4556 2324 4564
rect 2252 4536 2260 4544
rect 2284 4536 2292 4544
rect 2348 4536 2356 4544
rect 2156 4436 2164 4444
rect 2188 4436 2196 4444
rect 2076 4396 2084 4404
rect 2044 4356 2052 4364
rect 2060 4336 2068 4344
rect 2172 4356 2180 4364
rect 2188 4336 2196 4344
rect 2220 4376 2228 4384
rect 2252 4396 2260 4404
rect 2236 4356 2244 4364
rect 2380 4616 2388 4624
rect 2300 4516 2308 4524
rect 2364 4516 2372 4524
rect 2460 4596 2468 4604
rect 2540 4676 2548 4684
rect 2492 4476 2500 4484
rect 2444 4436 2452 4444
rect 2348 4416 2356 4424
rect 2380 4416 2388 4424
rect 2364 4376 2372 4384
rect 2396 4376 2404 4384
rect 2348 4356 2356 4364
rect 2268 4316 2276 4324
rect 2332 4316 2340 4324
rect 2012 4256 2020 4264
rect 1980 4096 1988 4104
rect 1884 3976 1892 3984
rect 1820 3916 1828 3924
rect 1948 3916 1956 3924
rect 1996 3936 2004 3944
rect 1996 3916 2004 3924
rect 2140 4296 2148 4304
rect 2204 4296 2212 4304
rect 2236 4296 2244 4304
rect 2204 4276 2212 4284
rect 2156 4256 2164 4264
rect 2028 4056 2036 4064
rect 2060 4056 2068 4064
rect 2044 4036 2052 4044
rect 2028 4016 2036 4024
rect 1692 3896 1700 3904
rect 1900 3896 1908 3904
rect 1932 3896 1940 3904
rect 1980 3896 1988 3904
rect 2012 3896 2020 3904
rect 1564 3856 1572 3864
rect 1468 3796 1476 3804
rect 1324 3756 1332 3764
rect 1340 3736 1348 3744
rect 1228 3696 1236 3704
rect 1276 3696 1284 3704
rect 1260 3656 1268 3664
rect 1052 3616 1060 3624
rect 940 3556 948 3564
rect 1020 3556 1028 3564
rect 1116 3556 1124 3564
rect 1084 3516 1092 3524
rect 876 3496 884 3504
rect 892 3496 900 3504
rect 924 3496 932 3504
rect 972 3496 980 3504
rect 1004 3496 1012 3504
rect 940 3476 948 3484
rect 1052 3476 1060 3484
rect 860 3456 868 3464
rect 908 3456 916 3464
rect 876 3436 884 3444
rect 924 3376 932 3384
rect 844 3356 852 3364
rect 860 3296 868 3304
rect 876 3236 884 3244
rect 876 3136 884 3144
rect 876 3096 884 3104
rect 956 3456 964 3464
rect 972 3436 980 3444
rect 940 3276 948 3284
rect 940 3216 948 3224
rect 1068 3356 1076 3364
rect 1020 3336 1028 3344
rect 1116 3456 1124 3464
rect 1180 3536 1188 3544
rect 1164 3516 1172 3524
rect 1196 3516 1204 3524
rect 1164 3496 1172 3504
rect 1052 3316 1060 3324
rect 1068 3316 1076 3324
rect 1100 3316 1108 3324
rect 1020 3296 1028 3304
rect 1004 3276 1012 3284
rect 1020 3256 1028 3264
rect 1132 3316 1140 3324
rect 1148 3316 1156 3324
rect 1084 3276 1092 3284
rect 1148 3276 1156 3284
rect 1180 3276 1188 3284
rect 972 3176 980 3184
rect 908 3136 916 3144
rect 1036 3116 1044 3124
rect 908 3096 916 3104
rect 988 3096 996 3104
rect 1068 3096 1076 3104
rect 940 3076 948 3084
rect 972 3016 980 3024
rect 940 2976 948 2984
rect 892 2956 900 2964
rect 860 2916 868 2924
rect 796 2756 804 2764
rect 764 2716 772 2724
rect 812 2716 820 2724
rect 540 2676 548 2684
rect 716 2656 724 2664
rect 828 2656 836 2664
rect 572 2636 580 2644
rect 540 2516 548 2524
rect 588 2516 596 2524
rect 588 2496 596 2504
rect 524 2476 532 2484
rect 668 2556 676 2564
rect 700 2556 708 2564
rect 812 2636 820 2644
rect 892 2896 900 2904
rect 876 2796 884 2804
rect 860 2756 868 2764
rect 940 2916 948 2924
rect 908 2876 916 2884
rect 924 2796 932 2804
rect 892 2716 900 2724
rect 844 2636 852 2644
rect 860 2636 868 2644
rect 828 2576 836 2584
rect 636 2516 644 2524
rect 764 2516 772 2524
rect 828 2516 836 2524
rect 684 2476 692 2484
rect 604 2436 612 2444
rect 524 2376 532 2384
rect 492 2356 500 2364
rect 460 2316 468 2324
rect 572 2336 580 2344
rect 620 2336 628 2344
rect 668 2356 676 2364
rect 540 2316 548 2324
rect 652 2316 660 2324
rect 764 2336 772 2344
rect 332 2296 340 2304
rect 364 2296 372 2304
rect 620 2296 628 2304
rect 716 2296 724 2304
rect 764 2296 772 2304
rect 428 2276 436 2284
rect 524 2276 532 2284
rect 460 2256 468 2264
rect 316 2136 324 2144
rect 252 2116 260 2124
rect 300 2116 308 2124
rect 284 2096 292 2104
rect 204 2076 212 2084
rect 172 1856 180 1864
rect 156 1836 164 1844
rect 204 1896 212 1904
rect 188 1816 196 1824
rect 252 1836 260 1844
rect 204 1796 212 1804
rect 316 2076 324 2084
rect 492 2256 500 2264
rect 572 2276 580 2284
rect 940 2776 948 2784
rect 1020 3076 1028 3084
rect 1004 2956 1012 2964
rect 1148 3156 1156 3164
rect 1116 3116 1124 3124
rect 1148 3096 1156 3104
rect 1164 3096 1172 3104
rect 1100 3076 1108 3084
rect 1148 3036 1156 3044
rect 1084 3016 1092 3024
rect 1116 3016 1124 3024
rect 1020 2936 1028 2944
rect 988 2896 996 2904
rect 1004 2876 1012 2884
rect 988 2816 996 2824
rect 1052 2916 1060 2924
rect 1084 2916 1092 2924
rect 1084 2876 1092 2884
rect 1100 2876 1108 2884
rect 1052 2836 1060 2844
rect 1100 2796 1108 2804
rect 1148 2936 1156 2944
rect 1036 2776 1044 2784
rect 1020 2756 1028 2764
rect 1004 2696 1012 2704
rect 956 2676 964 2684
rect 1020 2676 1028 2684
rect 908 2656 916 2664
rect 892 2496 900 2504
rect 1004 2656 1012 2664
rect 972 2636 980 2644
rect 956 2596 964 2604
rect 1068 2676 1076 2684
rect 1084 2636 1092 2644
rect 1084 2556 1092 2564
rect 1212 3456 1220 3464
rect 1212 3376 1220 3384
rect 1228 3356 1236 3364
rect 1212 3336 1220 3344
rect 1276 3556 1284 3564
rect 1260 3496 1268 3504
rect 1292 3496 1300 3504
rect 1276 3476 1284 3484
rect 1292 3436 1300 3444
rect 1324 3576 1332 3584
rect 1308 3356 1316 3364
rect 1308 3316 1316 3324
rect 1372 3696 1380 3704
rect 1500 3696 1508 3704
rect 1356 3636 1364 3644
rect 1388 3676 1396 3684
rect 1564 3696 1572 3704
rect 1724 3856 1732 3864
rect 1836 3856 1844 3864
rect 1692 3816 1700 3824
rect 1676 3776 1684 3784
rect 1724 3776 1732 3784
rect 1724 3716 1732 3724
rect 1644 3696 1652 3704
rect 1628 3676 1636 3684
rect 1660 3676 1668 3684
rect 1388 3656 1396 3664
rect 1516 3656 1524 3664
rect 1580 3656 1588 3664
rect 1372 3556 1380 3564
rect 1372 3536 1380 3544
rect 1468 3636 1476 3644
rect 1596 3636 1604 3644
rect 1411 3606 1419 3614
rect 1421 3606 1429 3614
rect 1431 3606 1439 3614
rect 1441 3606 1449 3614
rect 1451 3606 1459 3614
rect 1461 3606 1469 3614
rect 1452 3576 1460 3584
rect 1404 3556 1412 3564
rect 1388 3496 1396 3504
rect 1340 3476 1348 3484
rect 1388 3476 1396 3484
rect 1340 3456 1348 3464
rect 1356 3336 1364 3344
rect 1580 3616 1588 3624
rect 1548 3536 1556 3544
rect 1580 3536 1588 3544
rect 1516 3516 1524 3524
rect 1548 3516 1556 3524
rect 1484 3496 1492 3504
rect 1516 3496 1524 3504
rect 1484 3356 1492 3364
rect 1388 3316 1396 3324
rect 1500 3336 1508 3344
rect 1356 3296 1364 3304
rect 1324 3276 1332 3284
rect 1276 3236 1284 3244
rect 1244 3156 1252 3164
rect 1196 3116 1204 3124
rect 1212 3080 1220 3084
rect 1212 3076 1220 3080
rect 1196 2996 1204 3004
rect 1196 2976 1204 2984
rect 1228 2956 1236 2964
rect 1212 2936 1220 2944
rect 1196 2916 1204 2924
rect 1196 2876 1204 2884
rect 1148 2696 1156 2704
rect 1180 2696 1188 2704
rect 1164 2676 1172 2684
rect 1196 2676 1204 2684
rect 1148 2636 1156 2644
rect 1180 2636 1188 2644
rect 1164 2556 1172 2564
rect 924 2516 932 2524
rect 1052 2516 1060 2524
rect 1132 2516 1140 2524
rect 1180 2516 1188 2524
rect 908 2336 916 2344
rect 828 2296 836 2304
rect 876 2296 884 2304
rect 908 2296 916 2304
rect 732 2276 740 2284
rect 764 2276 772 2284
rect 780 2276 788 2284
rect 844 2276 852 2284
rect 876 2256 884 2264
rect 860 2236 868 2244
rect 492 2176 500 2184
rect 444 2136 452 2144
rect 380 2116 388 2124
rect 428 2116 436 2124
rect 396 2096 404 2104
rect 348 2036 356 2044
rect 348 1996 356 2004
rect 476 2116 484 2124
rect 652 2156 660 2164
rect 844 2216 852 2224
rect 684 2136 692 2144
rect 748 2136 756 2144
rect 828 2136 836 2144
rect 508 2116 516 2124
rect 540 2116 548 2124
rect 332 1916 340 1924
rect 428 1916 436 1924
rect 300 1876 308 1884
rect 188 1756 196 1764
rect 236 1756 244 1764
rect 60 1716 68 1724
rect 92 1716 100 1724
rect 60 1696 68 1704
rect 108 1696 116 1704
rect 28 1656 36 1664
rect 172 1736 180 1744
rect 204 1716 212 1724
rect 220 1716 228 1724
rect 156 1676 164 1684
rect 236 1676 244 1684
rect 316 1856 324 1864
rect 428 1856 436 1864
rect 540 2076 548 2084
rect 524 2056 532 2064
rect 556 2056 564 2064
rect 796 2116 804 2124
rect 620 2096 628 2104
rect 588 2036 596 2044
rect 668 2076 676 2084
rect 700 2076 708 2084
rect 908 2236 916 2244
rect 892 2136 900 2144
rect 972 2276 980 2284
rect 956 2216 964 2224
rect 940 2136 948 2144
rect 924 2096 932 2104
rect 812 2076 820 2084
rect 876 2076 884 2084
rect 924 2076 932 2084
rect 732 2056 740 2064
rect 732 2036 740 2044
rect 700 1976 708 1984
rect 508 1936 516 1944
rect 396 1816 404 1824
rect 444 1816 452 1824
rect 332 1796 340 1804
rect 428 1756 436 1764
rect 412 1716 420 1724
rect 428 1696 436 1704
rect 316 1676 324 1684
rect 492 1916 500 1924
rect 492 1876 500 1884
rect 668 1936 676 1944
rect 684 1916 692 1924
rect 620 1896 628 1904
rect 716 1896 724 1904
rect 684 1876 692 1884
rect 716 1876 724 1884
rect 636 1856 644 1864
rect 572 1776 580 1784
rect 476 1756 484 1764
rect 476 1736 484 1744
rect 572 1736 580 1744
rect 636 1736 644 1744
rect 540 1716 548 1724
rect 556 1716 564 1724
rect 268 1656 276 1664
rect 284 1656 292 1664
rect 460 1656 468 1664
rect 364 1556 372 1564
rect 412 1536 420 1544
rect 284 1496 292 1504
rect 348 1496 356 1504
rect 396 1496 404 1504
rect 44 1456 52 1464
rect 76 1456 84 1464
rect 172 1456 180 1464
rect 188 1456 196 1464
rect 300 1476 308 1484
rect 252 1456 260 1464
rect 140 1436 148 1444
rect 204 1436 212 1444
rect 76 1356 84 1364
rect 92 1356 100 1364
rect 140 1356 148 1364
rect 204 1356 212 1364
rect 220 1356 228 1364
rect 204 1336 212 1344
rect 124 1316 132 1324
rect 60 1276 68 1284
rect 92 1276 100 1284
rect 172 1256 180 1264
rect 172 1136 180 1144
rect 220 1316 228 1324
rect 236 1316 244 1324
rect 188 1116 196 1124
rect 12 1096 20 1104
rect 220 1096 228 1104
rect 60 1056 68 1064
rect 108 1036 116 1044
rect 156 1036 164 1044
rect 236 1036 244 1044
rect 316 1436 324 1444
rect 540 1496 548 1504
rect 620 1716 628 1724
rect 668 1716 676 1724
rect 716 1816 724 1824
rect 700 1776 708 1784
rect 780 1976 788 1984
rect 780 1956 788 1964
rect 764 1916 772 1924
rect 748 1856 756 1864
rect 1004 2376 1012 2384
rect 1196 2496 1204 2504
rect 1036 2356 1044 2364
rect 1020 2316 1028 2324
rect 1020 2236 1028 2244
rect 988 2176 996 2184
rect 1004 2136 1012 2144
rect 988 2076 996 2084
rect 940 2056 948 2064
rect 972 2056 980 2064
rect 956 1936 964 1944
rect 844 1880 852 1884
rect 844 1876 852 1880
rect 860 1856 868 1864
rect 700 1736 708 1744
rect 684 1576 692 1584
rect 636 1516 644 1524
rect 684 1516 692 1524
rect 572 1496 580 1504
rect 700 1496 708 1504
rect 492 1476 500 1484
rect 540 1476 548 1484
rect 572 1476 580 1484
rect 444 1456 452 1464
rect 492 1456 500 1464
rect 428 1436 436 1444
rect 460 1436 468 1444
rect 364 1376 372 1384
rect 300 1356 308 1364
rect 316 1356 324 1364
rect 556 1456 564 1464
rect 652 1436 660 1444
rect 556 1396 564 1404
rect 604 1396 612 1404
rect 332 1336 340 1344
rect 508 1336 516 1344
rect 364 1316 372 1324
rect 460 1316 468 1324
rect 492 1316 500 1324
rect 668 1396 676 1404
rect 908 1876 916 1884
rect 956 1916 964 1924
rect 1020 1936 1028 1944
rect 1004 1916 1012 1924
rect 972 1896 980 1904
rect 924 1856 932 1864
rect 972 1856 980 1864
rect 1004 1896 1012 1904
rect 1052 2276 1060 2284
rect 1180 2416 1188 2424
rect 1084 2376 1092 2384
rect 1116 2336 1124 2344
rect 1164 2316 1172 2324
rect 1132 2296 1140 2304
rect 1276 3096 1284 3104
rect 1276 3056 1284 3064
rect 1260 2956 1268 2964
rect 1372 3196 1380 3204
rect 1468 3256 1476 3264
rect 1516 3216 1524 3224
rect 1411 3206 1419 3214
rect 1421 3206 1429 3214
rect 1431 3206 1439 3214
rect 1441 3206 1449 3214
rect 1451 3206 1459 3214
rect 1461 3206 1469 3214
rect 1628 3576 1636 3584
rect 1628 3516 1636 3524
rect 1628 3376 1636 3384
rect 1596 3356 1604 3364
rect 1676 3596 1684 3604
rect 1740 3616 1748 3624
rect 1724 3496 1732 3504
rect 1708 3476 1716 3484
rect 1708 3396 1716 3404
rect 1708 3376 1716 3384
rect 1676 3316 1684 3324
rect 1660 3296 1668 3304
rect 1580 3276 1588 3284
rect 1612 3256 1620 3264
rect 1580 3236 1588 3244
rect 1532 3196 1540 3204
rect 1644 3216 1652 3224
rect 1948 3796 1956 3804
rect 1996 3796 2004 3804
rect 1836 3756 1844 3764
rect 1980 3756 1988 3764
rect 1820 3716 1828 3724
rect 2060 3936 2068 3944
rect 2044 3816 2052 3824
rect 1916 3736 1924 3744
rect 2012 3736 2020 3744
rect 1884 3716 1892 3724
rect 1996 3716 2004 3724
rect 1804 3576 1812 3584
rect 1772 3536 1780 3544
rect 1804 3536 1812 3544
rect 1756 3456 1764 3464
rect 1820 3376 1828 3384
rect 1820 3336 1828 3344
rect 1788 3316 1796 3324
rect 1740 3236 1748 3244
rect 1804 3256 1812 3264
rect 1772 3216 1780 3224
rect 1708 3196 1716 3204
rect 1724 3196 1732 3204
rect 1516 3176 1524 3184
rect 1612 3176 1620 3184
rect 1564 3156 1572 3164
rect 1500 3136 1508 3144
rect 1356 3116 1364 3124
rect 1276 2916 1284 2924
rect 1308 2916 1316 2924
rect 1244 2796 1252 2804
rect 1244 2636 1252 2644
rect 1244 2616 1252 2624
rect 1228 2456 1236 2464
rect 1196 2376 1204 2384
rect 1212 2376 1220 2384
rect 1100 2236 1108 2244
rect 1068 2176 1076 2184
rect 1068 2136 1076 2144
rect 1052 2076 1060 2084
rect 1132 2136 1140 2144
rect 1244 2396 1252 2404
rect 1244 2376 1252 2384
rect 1244 2356 1252 2364
rect 1228 2316 1236 2324
rect 1212 2256 1220 2264
rect 1244 2096 1252 2104
rect 1116 2076 1124 2084
rect 1292 2796 1300 2804
rect 1420 3076 1428 3084
rect 1516 3096 1524 3104
rect 1500 3056 1508 3064
rect 1532 3056 1540 3064
rect 1516 3036 1524 3044
rect 1500 3016 1508 3024
rect 1356 2996 1364 3004
rect 1356 2956 1364 2964
rect 1372 2956 1380 2964
rect 1276 2676 1284 2684
rect 1340 2756 1348 2764
rect 1324 2656 1332 2664
rect 1308 2636 1316 2644
rect 1292 2556 1300 2564
rect 1324 2556 1332 2564
rect 1276 2536 1284 2544
rect 1308 2536 1316 2544
rect 1308 2496 1316 2504
rect 1276 2296 1284 2304
rect 1308 2296 1316 2304
rect 1292 2256 1300 2264
rect 1308 2236 1316 2244
rect 1276 2156 1284 2164
rect 1260 2056 1268 2064
rect 1132 2016 1140 2024
rect 1116 1936 1124 1944
rect 1196 1936 1204 1944
rect 1212 1936 1220 1944
rect 1116 1916 1124 1924
rect 1164 1916 1172 1924
rect 1308 2116 1316 2124
rect 1308 2056 1316 2064
rect 1292 1996 1300 2004
rect 1276 1956 1284 1964
rect 1260 1896 1268 1904
rect 1052 1876 1060 1884
rect 1084 1876 1092 1884
rect 1340 2516 1348 2524
rect 1340 2296 1348 2304
rect 1340 2276 1348 2284
rect 1340 2256 1348 2264
rect 1468 2936 1476 2944
rect 1388 2916 1396 2924
rect 1372 2876 1380 2884
rect 1372 2776 1380 2784
rect 1411 2806 1419 2814
rect 1421 2806 1429 2814
rect 1431 2806 1439 2814
rect 1441 2806 1449 2814
rect 1451 2806 1459 2814
rect 1461 2806 1469 2814
rect 1596 3136 1604 3144
rect 1580 3096 1588 3104
rect 1580 2996 1588 3004
rect 1564 2936 1572 2944
rect 1900 3696 1908 3704
rect 1868 3576 1876 3584
rect 1884 3576 1892 3584
rect 1900 3556 1908 3564
rect 1884 3516 1892 3524
rect 2044 3516 2052 3524
rect 1948 3496 1956 3504
rect 2076 3516 2084 3524
rect 2076 3496 2084 3504
rect 1948 3456 1956 3464
rect 2012 3416 2020 3424
rect 1916 3396 1924 3404
rect 1884 3376 1892 3384
rect 1932 3356 1940 3364
rect 2012 3336 2020 3344
rect 1868 3296 1876 3304
rect 1916 3296 1924 3304
rect 1836 3276 1844 3284
rect 1836 3196 1844 3204
rect 2076 3376 2084 3384
rect 2108 4156 2116 4164
rect 2188 4136 2196 4144
rect 2124 4116 2132 4124
rect 2108 3956 2116 3964
rect 2188 3896 2196 3904
rect 2252 4196 2260 4204
rect 2380 4316 2388 4324
rect 2396 4316 2404 4324
rect 2780 5216 2788 5224
rect 2780 5196 2788 5204
rect 2796 5156 2804 5164
rect 2780 5016 2788 5024
rect 2732 4956 2740 4964
rect 2940 5276 2948 5284
rect 2988 5216 2996 5224
rect 2924 5136 2932 5144
rect 2844 5096 2852 5104
rect 2892 5096 2900 5104
rect 2812 5076 2820 5084
rect 2828 4956 2836 4964
rect 2716 4916 2724 4924
rect 2604 4856 2612 4864
rect 2620 4856 2628 4864
rect 2572 4836 2580 4844
rect 2604 4816 2612 4824
rect 2780 4896 2788 4904
rect 2700 4796 2708 4804
rect 2700 4756 2708 4764
rect 2668 4736 2676 4744
rect 2572 4716 2580 4724
rect 2556 4596 2564 4604
rect 2620 4616 2628 4624
rect 2588 4576 2596 4584
rect 2540 4556 2548 4564
rect 2540 4536 2548 4544
rect 2588 4536 2596 4544
rect 2652 4676 2660 4684
rect 2652 4656 2660 4664
rect 2684 4656 2692 4664
rect 2732 4676 2740 4684
rect 2716 4656 2724 4664
rect 2732 4616 2740 4624
rect 2684 4596 2692 4604
rect 2668 4576 2676 4584
rect 2876 5076 2884 5084
rect 2892 5016 2900 5024
rect 2915 5006 2923 5014
rect 2925 5006 2933 5014
rect 2935 5006 2943 5014
rect 2945 5006 2953 5014
rect 2955 5006 2963 5014
rect 2965 5006 2973 5014
rect 3436 5416 3444 5424
rect 3500 5416 3508 5424
rect 3436 5396 3444 5404
rect 3468 5396 3476 5404
rect 3564 5396 3572 5404
rect 3356 5376 3364 5384
rect 3068 5356 3076 5364
rect 3100 5336 3108 5344
rect 3212 5336 3220 5344
rect 3340 5336 3348 5344
rect 3132 5156 3140 5164
rect 3324 5296 3332 5304
rect 3404 5356 3412 5364
rect 3420 5336 3428 5344
rect 3452 5376 3460 5384
rect 3468 5336 3476 5344
rect 3548 5336 3556 5344
rect 3372 5296 3380 5304
rect 3500 5316 3508 5324
rect 3564 5316 3572 5324
rect 3436 5276 3444 5284
rect 3452 5276 3460 5284
rect 3260 5136 3268 5144
rect 3052 5116 3060 5124
rect 3212 5116 3220 5124
rect 3036 4996 3044 5004
rect 3100 4996 3108 5004
rect 2892 4936 2900 4944
rect 3052 4936 3060 4944
rect 2860 4776 2868 4784
rect 2844 4736 2852 4744
rect 2764 4696 2772 4704
rect 2828 4696 2836 4704
rect 2876 4696 2884 4704
rect 2780 4676 2788 4684
rect 2876 4596 2884 4604
rect 2764 4576 2772 4584
rect 2780 4576 2788 4584
rect 2748 4556 2756 4564
rect 2860 4556 2868 4564
rect 2572 4516 2580 4524
rect 2764 4536 2772 4544
rect 2828 4536 2836 4544
rect 2636 4516 2644 4524
rect 2748 4516 2756 4524
rect 2796 4516 2804 4524
rect 2716 4496 2724 4504
rect 2620 4456 2628 4464
rect 2604 4436 2612 4444
rect 2556 4396 2564 4404
rect 2476 4316 2484 4324
rect 2540 4316 2548 4324
rect 2396 4296 2404 4304
rect 2428 4296 2436 4304
rect 2364 4276 2372 4284
rect 2316 4256 2324 4264
rect 2348 4256 2356 4264
rect 2220 4176 2228 4184
rect 2252 4176 2260 4184
rect 2268 4176 2276 4184
rect 2236 4156 2244 4164
rect 2316 4136 2324 4144
rect 2236 4116 2244 4124
rect 2284 4116 2292 4124
rect 2348 4116 2356 4124
rect 2460 4276 2468 4284
rect 2508 4276 2516 4284
rect 2428 4236 2436 4244
rect 2460 4236 2468 4244
rect 2412 4216 2420 4224
rect 2428 4136 2436 4144
rect 2412 4116 2420 4124
rect 2380 4076 2388 4084
rect 2284 3936 2292 3944
rect 2364 3936 2372 3944
rect 2236 3896 2244 3904
rect 2524 4236 2532 4244
rect 2476 4216 2484 4224
rect 2476 4176 2484 4184
rect 2460 4156 2468 4164
rect 2476 4076 2484 4084
rect 2476 3896 2484 3904
rect 2524 4156 2532 4164
rect 2700 4396 2708 4404
rect 2572 4296 2580 4304
rect 2604 4296 2612 4304
rect 2588 4236 2596 4244
rect 2572 4196 2580 4204
rect 2684 4316 2692 4324
rect 2652 4296 2660 4304
rect 2668 4256 2676 4264
rect 2732 4316 2740 4324
rect 2748 4256 2756 4264
rect 2732 4196 2740 4204
rect 2700 4176 2708 4184
rect 2620 4156 2628 4164
rect 2556 4136 2564 4144
rect 2572 4136 2580 4144
rect 2636 4136 2644 4144
rect 2540 4116 2548 4124
rect 2508 3996 2516 4004
rect 2508 3936 2516 3944
rect 2572 4076 2580 4084
rect 2604 4056 2612 4064
rect 2620 3916 2628 3924
rect 2556 3896 2564 3904
rect 2316 3876 2324 3884
rect 2380 3876 2388 3884
rect 2604 3876 2612 3884
rect 2140 3856 2148 3864
rect 2140 3736 2148 3744
rect 2284 3856 2292 3864
rect 2620 3836 2628 3844
rect 2204 3796 2212 3804
rect 2220 3796 2228 3804
rect 2268 3796 2276 3804
rect 2316 3796 2324 3804
rect 2204 3736 2212 3744
rect 2156 3716 2164 3724
rect 2124 3696 2132 3704
rect 2108 3656 2116 3664
rect 2204 3656 2212 3664
rect 2092 3316 2100 3324
rect 1996 3296 2004 3304
rect 1964 3276 1972 3284
rect 2012 3276 2020 3284
rect 2028 3276 2036 3284
rect 2060 3276 2068 3284
rect 1948 3256 1956 3264
rect 1964 3256 1972 3264
rect 1932 3196 1940 3204
rect 1660 3136 1668 3144
rect 1724 3136 1732 3144
rect 1788 3136 1796 3144
rect 1852 3136 1860 3144
rect 1692 3096 1700 3104
rect 1644 3036 1652 3044
rect 1644 2976 1652 2984
rect 1660 2956 1668 2964
rect 1676 2936 1684 2944
rect 1708 3036 1716 3044
rect 1772 3036 1780 3044
rect 1724 3016 1732 3024
rect 1708 2956 1716 2964
rect 1740 2936 1748 2944
rect 1548 2916 1556 2924
rect 1644 2916 1652 2924
rect 1740 2916 1748 2924
rect 1612 2876 1620 2884
rect 1596 2816 1604 2824
rect 1532 2796 1540 2804
rect 1500 2736 1508 2744
rect 1388 2696 1396 2704
rect 1388 2516 1396 2524
rect 1420 2556 1428 2564
rect 1436 2496 1444 2504
rect 1420 2456 1428 2464
rect 1436 2456 1444 2464
rect 1411 2406 1419 2414
rect 1421 2406 1429 2414
rect 1431 2406 1439 2414
rect 1441 2406 1449 2414
rect 1451 2406 1459 2414
rect 1461 2406 1469 2414
rect 1420 2316 1428 2324
rect 1468 2296 1476 2304
rect 1452 2276 1460 2284
rect 1468 2216 1476 2224
rect 1340 2156 1348 2164
rect 1404 2156 1412 2164
rect 1356 2116 1364 2124
rect 1404 2096 1412 2104
rect 1436 2056 1444 2064
rect 1324 2036 1332 2044
rect 1324 1976 1332 1984
rect 1411 2006 1419 2014
rect 1421 2006 1429 2014
rect 1431 2006 1439 2014
rect 1441 2006 1449 2014
rect 1451 2006 1459 2014
rect 1461 2006 1469 2014
rect 1372 1996 1380 2004
rect 1356 1976 1364 1984
rect 1372 1976 1380 1984
rect 1308 1956 1316 1964
rect 1340 1956 1348 1964
rect 1324 1936 1332 1944
rect 1308 1896 1316 1904
rect 1340 1896 1348 1904
rect 1036 1856 1044 1864
rect 1068 1856 1076 1864
rect 988 1836 996 1844
rect 940 1776 948 1784
rect 1116 1776 1124 1784
rect 1052 1756 1060 1764
rect 1084 1756 1092 1764
rect 780 1716 788 1724
rect 780 1576 788 1584
rect 748 1536 756 1544
rect 764 1496 772 1504
rect 828 1696 836 1704
rect 748 1456 756 1464
rect 812 1476 820 1484
rect 844 1516 852 1524
rect 908 1736 916 1744
rect 940 1736 948 1744
rect 876 1516 884 1524
rect 860 1476 868 1484
rect 876 1476 884 1484
rect 828 1456 836 1464
rect 844 1456 852 1464
rect 796 1416 804 1424
rect 732 1376 740 1384
rect 636 1356 644 1364
rect 700 1356 708 1364
rect 860 1396 868 1404
rect 1004 1716 1012 1724
rect 940 1656 948 1664
rect 924 1536 932 1544
rect 924 1516 932 1524
rect 908 1476 916 1484
rect 972 1476 980 1484
rect 972 1456 980 1464
rect 748 1336 756 1344
rect 796 1336 804 1344
rect 844 1336 852 1344
rect 908 1336 916 1344
rect 540 1296 548 1304
rect 620 1296 628 1304
rect 284 1276 292 1284
rect 364 1276 372 1284
rect 588 1276 596 1284
rect 604 1276 612 1284
rect 668 1276 676 1284
rect 300 1256 308 1264
rect 284 1076 292 1084
rect 268 1056 276 1064
rect 284 1036 292 1044
rect 732 1136 740 1144
rect 492 1116 500 1124
rect 668 1116 676 1124
rect 780 1316 788 1324
rect 892 1316 900 1324
rect 940 1316 948 1324
rect 828 1276 836 1284
rect 796 1216 804 1224
rect 844 1136 852 1144
rect 1084 1696 1092 1704
rect 1068 1576 1076 1584
rect 1100 1536 1108 1544
rect 1068 1516 1076 1524
rect 1036 1476 1044 1484
rect 1084 1496 1092 1504
rect 1068 1456 1076 1464
rect 1100 1436 1108 1444
rect 1004 1356 1012 1364
rect 1212 1856 1220 1864
rect 1244 1856 1252 1864
rect 1228 1836 1236 1844
rect 1148 1756 1156 1764
rect 1180 1736 1188 1744
rect 1148 1716 1156 1724
rect 1132 1696 1140 1704
rect 1260 1756 1268 1764
rect 1260 1576 1268 1584
rect 1148 1536 1156 1544
rect 1228 1476 1236 1484
rect 1164 1436 1172 1444
rect 1180 1436 1188 1444
rect 1212 1436 1220 1444
rect 1260 1436 1268 1444
rect 1212 1376 1220 1384
rect 1148 1356 1156 1364
rect 1020 1196 1028 1204
rect 1132 1316 1140 1324
rect 1212 1336 1220 1344
rect 1260 1316 1268 1324
rect 1180 1256 1188 1264
rect 1052 1156 1060 1164
rect 956 1136 964 1144
rect 972 1136 980 1144
rect 956 1116 964 1124
rect 316 1096 324 1104
rect 364 1096 372 1104
rect 444 1096 452 1104
rect 652 1096 660 1104
rect 684 1096 692 1104
rect 908 1096 916 1104
rect 332 1056 340 1064
rect 316 1036 324 1044
rect 220 996 228 1004
rect 124 976 132 984
rect 156 976 164 984
rect 284 936 292 944
rect 12 896 20 904
rect 44 876 52 884
rect 12 856 20 864
rect 60 856 68 864
rect 108 716 116 724
rect 236 916 244 924
rect 156 716 164 724
rect 60 676 68 684
rect 140 676 148 684
rect 156 676 164 684
rect 76 656 84 664
rect 156 656 164 664
rect 188 676 196 684
rect 76 636 84 644
rect 108 576 116 584
rect 28 556 36 564
rect 60 556 68 564
rect 44 536 52 544
rect 188 536 196 544
rect 44 516 52 524
rect 252 636 260 644
rect 236 616 244 624
rect 236 576 244 584
rect 428 1076 436 1084
rect 396 1056 404 1064
rect 364 1016 372 1024
rect 364 936 372 944
rect 444 916 452 924
rect 332 896 340 904
rect 364 896 372 904
rect 396 876 404 884
rect 316 736 324 744
rect 508 1056 516 1064
rect 540 1056 548 1064
rect 556 1056 564 1064
rect 572 1056 580 1064
rect 636 1056 644 1064
rect 508 1036 516 1044
rect 476 956 484 964
rect 492 916 500 924
rect 460 856 468 864
rect 492 856 500 864
rect 364 696 372 704
rect 412 696 420 704
rect 460 716 468 724
rect 284 676 292 684
rect 300 656 308 664
rect 364 656 372 664
rect 396 636 404 644
rect 284 556 292 564
rect 380 556 388 564
rect 348 536 356 544
rect 364 536 372 544
rect 44 496 52 504
rect 140 496 148 504
rect 204 496 212 504
rect 268 516 276 524
rect 236 476 244 484
rect 108 296 116 304
rect 12 276 20 284
rect 60 236 68 244
rect 108 236 116 244
rect 124 236 132 244
rect 300 496 308 504
rect 332 496 340 504
rect 380 496 388 504
rect 460 676 468 684
rect 476 676 484 684
rect 476 636 484 644
rect 524 976 532 984
rect 556 1016 564 1024
rect 524 956 532 964
rect 588 956 596 964
rect 620 956 628 964
rect 652 956 660 964
rect 684 956 692 964
rect 652 936 660 944
rect 572 916 580 924
rect 668 916 676 924
rect 556 896 564 904
rect 716 936 724 944
rect 732 916 740 924
rect 540 736 548 744
rect 524 716 532 724
rect 540 696 548 704
rect 572 736 580 744
rect 572 696 580 704
rect 668 696 676 704
rect 684 696 692 704
rect 780 1056 788 1064
rect 860 1076 868 1084
rect 828 1036 836 1044
rect 764 1016 772 1024
rect 796 1016 804 1024
rect 1020 1116 1028 1124
rect 1068 1096 1076 1104
rect 1084 1096 1092 1104
rect 1148 1096 1156 1104
rect 1052 1076 1060 1084
rect 796 996 804 1004
rect 876 996 884 1004
rect 812 976 820 984
rect 876 976 884 984
rect 780 956 788 964
rect 860 956 868 964
rect 892 956 900 964
rect 988 1056 996 1064
rect 972 1036 980 1044
rect 1052 1016 1060 1024
rect 1116 1076 1124 1084
rect 1084 1056 1092 1064
rect 1164 1036 1172 1044
rect 1100 1016 1108 1024
rect 860 876 868 884
rect 844 836 852 844
rect 812 716 820 724
rect 876 716 884 724
rect 412 536 420 544
rect 508 536 516 544
rect 412 496 420 504
rect 716 676 724 684
rect 940 956 948 964
rect 956 956 964 964
rect 1036 956 1044 964
rect 1100 996 1108 1004
rect 956 936 964 944
rect 1068 936 1076 944
rect 924 916 932 924
rect 1020 916 1028 924
rect 940 836 948 844
rect 924 796 932 804
rect 748 656 756 664
rect 780 656 788 664
rect 796 656 804 664
rect 700 596 708 604
rect 780 636 788 644
rect 556 556 564 564
rect 684 556 692 564
rect 700 556 708 564
rect 748 556 756 564
rect 908 676 916 684
rect 844 656 852 664
rect 812 636 820 644
rect 844 596 852 604
rect 860 556 868 564
rect 908 556 916 564
rect 620 536 628 544
rect 700 536 708 544
rect 588 516 596 524
rect 652 516 660 524
rect 876 516 884 524
rect 1020 756 1028 764
rect 956 716 964 724
rect 940 676 948 684
rect 956 676 964 684
rect 1004 676 1012 684
rect 940 556 948 564
rect 668 496 676 504
rect 716 496 724 504
rect 748 496 756 504
rect 844 496 852 504
rect 876 496 884 504
rect 396 336 404 344
rect 364 316 372 324
rect 428 316 436 324
rect 236 296 244 304
rect 284 296 292 304
rect 348 296 356 304
rect 204 276 212 284
rect 188 236 196 244
rect 204 236 212 244
rect 188 196 196 204
rect 140 176 148 184
rect 156 156 164 164
rect 12 136 20 144
rect 44 136 52 144
rect 92 136 100 144
rect 76 116 84 124
rect 124 116 132 124
rect 252 256 260 264
rect 220 196 228 204
rect 220 176 228 184
rect 780 376 788 384
rect 748 356 756 364
rect 668 336 676 344
rect 572 316 580 324
rect 572 296 580 304
rect 604 296 612 304
rect 396 276 404 284
rect 460 276 468 284
rect 316 256 324 264
rect 300 236 308 244
rect 428 236 436 244
rect 332 196 340 204
rect 332 156 340 164
rect 348 156 356 164
rect 460 216 468 224
rect 524 256 532 264
rect 412 176 420 184
rect 508 176 516 184
rect 508 156 516 164
rect 588 276 596 284
rect 636 276 644 284
rect 652 276 660 284
rect 684 316 692 324
rect 700 276 708 284
rect 716 276 724 284
rect 652 236 660 244
rect 668 236 676 244
rect 604 196 612 204
rect 636 216 644 224
rect 620 176 628 184
rect 764 296 772 304
rect 844 336 852 344
rect 796 316 804 324
rect 844 316 852 324
rect 892 316 900 324
rect 972 656 980 664
rect 1036 716 1044 724
rect 1052 676 1060 684
rect 1036 656 1044 664
rect 1068 656 1076 664
rect 1084 656 1092 664
rect 988 576 996 584
rect 1004 536 1012 544
rect 1036 516 1044 524
rect 972 496 980 504
rect 1052 476 1060 484
rect 1116 956 1124 964
rect 1324 1876 1332 1884
rect 1388 1956 1396 1964
rect 1516 2496 1524 2504
rect 1564 2696 1572 2704
rect 1692 2896 1700 2904
rect 1820 3116 1828 3124
rect 1852 3116 1860 3124
rect 1804 3036 1812 3044
rect 1836 3036 1844 3044
rect 1820 2996 1828 3004
rect 1948 3156 1956 3164
rect 1884 3076 1892 3084
rect 1868 3036 1876 3044
rect 1868 2976 1876 2984
rect 1820 2916 1828 2924
rect 1772 2876 1780 2884
rect 1676 2776 1684 2784
rect 1724 2776 1732 2784
rect 1644 2756 1652 2764
rect 1660 2756 1668 2764
rect 1644 2696 1652 2704
rect 1548 2576 1556 2584
rect 1548 2556 1556 2564
rect 1564 2536 1572 2544
rect 1548 2496 1556 2504
rect 1532 2436 1540 2444
rect 1772 2776 1780 2784
rect 1708 2736 1716 2744
rect 1868 2756 1876 2764
rect 1804 2716 1812 2724
rect 1708 2696 1716 2704
rect 1756 2696 1764 2704
rect 1612 2576 1620 2584
rect 1628 2556 1636 2564
rect 1596 2536 1604 2544
rect 1628 2496 1636 2504
rect 1660 2656 1668 2664
rect 1580 2456 1588 2464
rect 1612 2436 1620 2444
rect 1516 2356 1524 2364
rect 1532 2336 1540 2344
rect 1548 2336 1556 2344
rect 1868 2676 1876 2684
rect 1788 2616 1796 2624
rect 1852 2636 1860 2644
rect 1820 2576 1828 2584
rect 1836 2576 1844 2584
rect 1724 2556 1732 2564
rect 1756 2556 1764 2564
rect 1868 2556 1876 2564
rect 1740 2536 1748 2544
rect 1852 2536 1860 2544
rect 1932 3056 1940 3064
rect 1964 3056 1972 3064
rect 1900 2976 1908 2984
rect 2012 3216 2020 3224
rect 2012 3076 2020 3084
rect 1980 3016 1988 3024
rect 1964 2956 1972 2964
rect 2076 3216 2084 3224
rect 2060 3096 2068 3104
rect 2012 2936 2020 2944
rect 2028 2936 2036 2944
rect 1980 2916 1988 2924
rect 2060 2916 2068 2924
rect 1948 2816 1956 2824
rect 1916 2776 1924 2784
rect 1948 2756 1956 2764
rect 1900 2536 1908 2544
rect 1580 2316 1588 2324
rect 1660 2316 1668 2324
rect 1532 2236 1540 2244
rect 1516 2116 1524 2124
rect 1516 2096 1524 2104
rect 1564 2076 1572 2084
rect 1564 2056 1572 2064
rect 1548 1976 1556 1984
rect 1596 2096 1604 2104
rect 1660 2276 1668 2284
rect 1628 2176 1636 2184
rect 1628 2076 1636 2084
rect 1612 2056 1620 2064
rect 1596 2016 1604 2024
rect 1564 1956 1572 1964
rect 1580 1956 1588 1964
rect 1612 1956 1620 1964
rect 1372 1896 1380 1904
rect 1356 1856 1364 1864
rect 1292 1796 1300 1804
rect 1356 1796 1364 1804
rect 1388 1796 1396 1804
rect 1308 1756 1316 1764
rect 1324 1756 1332 1764
rect 1340 1756 1348 1764
rect 1292 1696 1300 1704
rect 1500 1796 1508 1804
rect 1516 1796 1524 1804
rect 1644 2016 1652 2024
rect 1644 1916 1652 1924
rect 1628 1896 1636 1904
rect 1628 1776 1636 1784
rect 1404 1756 1412 1764
rect 1548 1736 1556 1744
rect 1516 1716 1524 1724
rect 1532 1716 1540 1724
rect 1356 1676 1364 1684
rect 1500 1676 1508 1684
rect 1484 1636 1492 1644
rect 1411 1606 1419 1614
rect 1421 1606 1429 1614
rect 1431 1606 1439 1614
rect 1441 1606 1449 1614
rect 1451 1606 1459 1614
rect 1461 1606 1469 1614
rect 1308 1496 1316 1504
rect 1292 1376 1300 1384
rect 1324 1476 1332 1484
rect 1340 1436 1348 1444
rect 1340 1396 1348 1404
rect 1324 1356 1332 1364
rect 1212 1236 1220 1244
rect 1244 1236 1252 1244
rect 1276 1236 1284 1244
rect 1212 1216 1220 1224
rect 1196 936 1204 944
rect 1228 1076 1236 1084
rect 1372 1336 1380 1344
rect 1372 1296 1380 1304
rect 1692 2336 1700 2344
rect 1740 2436 1748 2444
rect 1852 2516 1860 2524
rect 1884 2516 1892 2524
rect 1740 2376 1748 2384
rect 1756 2376 1764 2384
rect 1724 2276 1732 2284
rect 1788 2336 1796 2344
rect 1772 2276 1780 2284
rect 1740 2256 1748 2264
rect 1692 2116 1700 2124
rect 1676 2096 1684 2104
rect 1692 2096 1700 2104
rect 1676 2076 1684 2084
rect 1708 2076 1716 2084
rect 1708 2036 1716 2044
rect 1676 1956 1684 1964
rect 1724 1956 1732 1964
rect 1692 1896 1700 1904
rect 1692 1876 1700 1884
rect 1676 1716 1684 1724
rect 1580 1656 1588 1664
rect 1692 1676 1700 1684
rect 1740 1876 1748 1884
rect 1740 1756 1748 1764
rect 1884 2476 1892 2484
rect 1884 2396 1892 2404
rect 1932 2556 1940 2564
rect 2044 2856 2052 2864
rect 2012 2836 2020 2844
rect 1996 2656 2004 2664
rect 1948 2536 1956 2544
rect 1980 2556 1988 2564
rect 2060 2636 2068 2644
rect 2044 2616 2052 2624
rect 2028 2556 2036 2564
rect 2012 2536 2020 2544
rect 1916 2476 1924 2484
rect 1932 2356 1940 2364
rect 1900 2296 1908 2304
rect 1868 2276 1876 2284
rect 1900 2276 1908 2284
rect 1852 2256 1860 2264
rect 1964 2336 1972 2344
rect 2268 3776 2276 3784
rect 2252 3756 2260 3764
rect 2332 3736 2340 3744
rect 2412 3736 2420 3744
rect 2300 3716 2308 3724
rect 2348 3716 2356 3724
rect 2300 3556 2308 3564
rect 2252 3536 2260 3544
rect 2300 3516 2308 3524
rect 2236 3496 2244 3504
rect 2220 3456 2228 3464
rect 2364 3656 2372 3664
rect 2396 3656 2404 3664
rect 2364 3536 2372 3544
rect 2332 3496 2340 3504
rect 2364 3496 2372 3504
rect 2332 3476 2340 3484
rect 2348 3456 2356 3464
rect 2188 3436 2196 3444
rect 2300 3436 2308 3444
rect 2140 3296 2148 3304
rect 2108 3216 2116 3224
rect 2140 3196 2148 3204
rect 2156 3156 2164 3164
rect 2124 3136 2132 3144
rect 2156 3136 2164 3144
rect 2092 3116 2100 3124
rect 2108 3056 2116 3064
rect 2236 3416 2244 3424
rect 2188 3356 2196 3364
rect 2252 3356 2260 3364
rect 2236 3336 2244 3344
rect 2460 3816 2468 3824
rect 2444 3756 2452 3764
rect 2556 3736 2564 3744
rect 2492 3716 2500 3724
rect 2524 3716 2532 3724
rect 2652 4116 2660 4124
rect 2668 4016 2676 4024
rect 2796 4436 2804 4444
rect 2796 4376 2804 4384
rect 2780 4276 2788 4284
rect 2780 4216 2788 4224
rect 2764 4176 2772 4184
rect 2796 4176 2804 4184
rect 2924 4856 2932 4864
rect 2988 4836 2996 4844
rect 3052 4876 3060 4884
rect 3036 4796 3044 4804
rect 2988 4676 2996 4684
rect 3004 4656 3012 4664
rect 2988 4616 2996 4624
rect 2915 4606 2923 4614
rect 2925 4606 2933 4614
rect 2935 4606 2943 4614
rect 2945 4606 2953 4614
rect 2955 4606 2963 4614
rect 2965 4606 2973 4614
rect 2892 4516 2900 4524
rect 2924 4536 2932 4544
rect 2908 4436 2916 4444
rect 2892 4376 2900 4384
rect 2876 4316 2884 4324
rect 2892 4296 2900 4304
rect 3020 4556 3028 4564
rect 3004 4516 3012 4524
rect 3004 4496 3012 4504
rect 3084 4836 3092 4844
rect 3068 4696 3076 4704
rect 3084 4616 3092 4624
rect 3132 4876 3140 4884
rect 3244 5096 3252 5104
rect 3180 5056 3188 5064
rect 3228 5016 3236 5024
rect 3196 4916 3204 4924
rect 3244 4896 3252 4904
rect 3308 5116 3316 5124
rect 3276 4996 3284 5004
rect 3292 4956 3300 4964
rect 3276 4916 3284 4924
rect 3324 4916 3332 4924
rect 3164 4876 3172 4884
rect 3260 4876 3268 4884
rect 3164 4836 3172 4844
rect 3148 4696 3156 4704
rect 3132 4656 3140 4664
rect 3180 4656 3188 4664
rect 3068 4536 3076 4544
rect 3132 4536 3140 4544
rect 3036 4496 3044 4504
rect 3052 4496 3060 4504
rect 3052 4476 3060 4484
rect 3020 4376 3028 4384
rect 2988 4296 2996 4304
rect 2988 4236 2996 4244
rect 2915 4206 2923 4214
rect 2925 4206 2933 4214
rect 2935 4206 2943 4214
rect 2945 4206 2953 4214
rect 2955 4206 2963 4214
rect 2965 4206 2973 4214
rect 2908 4176 2916 4184
rect 2828 4156 2836 4164
rect 2860 4156 2868 4164
rect 2780 4136 2788 4144
rect 2828 4136 2836 4144
rect 2748 4116 2756 4124
rect 2812 4116 2820 4124
rect 2924 4156 2932 4164
rect 2764 4076 2772 4084
rect 2844 4076 2852 4084
rect 2732 4016 2740 4024
rect 2732 3996 2740 4004
rect 2700 3896 2708 3904
rect 2652 3876 2660 3884
rect 2716 3876 2724 3884
rect 2876 4016 2884 4024
rect 2844 3996 2852 4004
rect 2796 3916 2804 3924
rect 2764 3876 2772 3884
rect 2668 3796 2676 3804
rect 2636 3776 2644 3784
rect 2716 3736 2724 3744
rect 2780 3816 2788 3824
rect 2780 3796 2788 3804
rect 2748 3736 2756 3744
rect 2844 3896 2852 3904
rect 2988 4096 2996 4104
rect 2988 3956 2996 3964
rect 2860 3876 2868 3884
rect 2876 3876 2884 3884
rect 3004 3876 3012 3884
rect 2988 3856 2996 3864
rect 3004 3836 3012 3844
rect 2915 3806 2923 3814
rect 2925 3806 2933 3814
rect 2935 3806 2943 3814
rect 2945 3806 2953 3814
rect 2955 3806 2963 3814
rect 2965 3806 2973 3814
rect 2876 3796 2884 3804
rect 2876 3756 2884 3764
rect 2812 3736 2820 3744
rect 2908 3736 2916 3744
rect 2604 3716 2612 3724
rect 2620 3716 2628 3724
rect 2524 3556 2532 3564
rect 2460 3516 2468 3524
rect 2492 3516 2500 3524
rect 2492 3476 2500 3484
rect 2508 3456 2516 3464
rect 2476 3416 2484 3424
rect 2460 3376 2468 3384
rect 2284 3316 2292 3324
rect 2204 3276 2212 3284
rect 2140 2976 2148 2984
rect 2188 2976 2196 2984
rect 2108 2936 2116 2944
rect 2092 2816 2100 2824
rect 2108 2696 2116 2704
rect 2316 3216 2324 3224
rect 2300 3136 2308 3144
rect 2236 3116 2244 3124
rect 2396 3336 2404 3344
rect 2428 3336 2436 3344
rect 2348 3316 2356 3324
rect 2300 3116 2308 3124
rect 2332 3116 2340 3124
rect 2316 3096 2324 3104
rect 2332 3096 2340 3104
rect 2220 3056 2228 3064
rect 2284 3056 2292 3064
rect 2236 2936 2244 2944
rect 2300 2936 2308 2944
rect 2204 2856 2212 2864
rect 2284 2856 2292 2864
rect 2300 2856 2308 2864
rect 2140 2716 2148 2724
rect 2124 2596 2132 2604
rect 2092 2556 2100 2564
rect 2028 2476 2036 2484
rect 2012 2456 2020 2464
rect 1964 2316 1972 2324
rect 1788 2176 1796 2184
rect 1852 2176 1860 2184
rect 1900 2176 1908 2184
rect 1916 2176 1924 2184
rect 1772 2156 1780 2164
rect 1852 2096 1860 2104
rect 1868 2096 1876 2104
rect 1772 2076 1780 2084
rect 1804 2076 1812 2084
rect 1788 2036 1796 2044
rect 1932 2096 1940 2104
rect 1964 2096 1972 2104
rect 1852 2056 1860 2064
rect 1916 2056 1924 2064
rect 1916 2016 1924 2024
rect 1836 1976 1844 1984
rect 1900 1976 1908 1984
rect 1916 1976 1924 1984
rect 1852 1956 1860 1964
rect 1916 1956 1924 1964
rect 1788 1896 1796 1904
rect 1964 1936 1972 1944
rect 1996 2316 2004 2324
rect 2044 2316 2052 2324
rect 2044 2276 2052 2284
rect 2156 2596 2164 2604
rect 2220 2716 2228 2724
rect 2268 2696 2276 2704
rect 2204 2616 2212 2624
rect 2204 2576 2212 2584
rect 2380 3156 2388 3164
rect 2380 3076 2388 3084
rect 2428 3316 2436 3324
rect 2412 3296 2420 3304
rect 2444 3236 2452 3244
rect 2460 3236 2468 3244
rect 2444 3156 2452 3164
rect 2412 3136 2420 3144
rect 2556 3496 2564 3504
rect 2588 3496 2596 3504
rect 2636 3636 2644 3644
rect 2572 3476 2580 3484
rect 2572 3356 2580 3364
rect 2556 3316 2564 3324
rect 2508 3296 2516 3304
rect 2492 3256 2500 3264
rect 2492 3136 2500 3144
rect 2428 3116 2436 3124
rect 2476 3116 2484 3124
rect 2412 3096 2420 3104
rect 2476 3096 2484 3104
rect 2396 2996 2404 3004
rect 2396 2976 2404 2984
rect 2364 2896 2372 2904
rect 2396 2896 2404 2904
rect 2332 2836 2340 2844
rect 2428 2996 2436 3004
rect 2540 3156 2548 3164
rect 2556 3136 2564 3144
rect 2524 3116 2532 3124
rect 2540 3076 2548 3084
rect 2540 3056 2548 3064
rect 2508 3036 2516 3044
rect 2524 3036 2532 3044
rect 2556 2976 2564 2984
rect 2476 2896 2484 2904
rect 2476 2876 2484 2884
rect 2508 2876 2516 2884
rect 2412 2816 2420 2824
rect 2396 2716 2404 2724
rect 2444 2716 2452 2724
rect 2396 2656 2404 2664
rect 2476 2676 2484 2684
rect 2476 2656 2484 2664
rect 2460 2636 2468 2644
rect 2332 2616 2340 2624
rect 2284 2556 2292 2564
rect 2236 2516 2244 2524
rect 2204 2496 2212 2504
rect 2220 2496 2228 2504
rect 2236 2476 2244 2484
rect 2364 2596 2372 2604
rect 2396 2616 2404 2624
rect 2380 2536 2388 2544
rect 2204 2456 2212 2464
rect 2268 2456 2276 2464
rect 2124 2316 2132 2324
rect 2156 2336 2164 2344
rect 2092 2296 2100 2304
rect 2076 2176 2084 2184
rect 2108 2276 2116 2284
rect 2108 2176 2116 2184
rect 2028 2156 2036 2164
rect 2044 2136 2052 2144
rect 1996 2056 2004 2064
rect 2060 2056 2068 2064
rect 2028 2036 2036 2044
rect 2076 2036 2084 2044
rect 2108 1996 2116 2004
rect 2140 2276 2148 2284
rect 2140 2176 2148 2184
rect 2268 2336 2276 2344
rect 2300 2336 2308 2344
rect 2268 2316 2276 2324
rect 2268 2296 2276 2304
rect 2332 2496 2340 2504
rect 2428 2556 2436 2564
rect 2540 2856 2548 2864
rect 2556 2716 2564 2724
rect 2620 3356 2628 3364
rect 2732 3536 2740 3544
rect 2684 3496 2692 3504
rect 2732 3476 2740 3484
rect 2716 3356 2724 3364
rect 2636 3336 2644 3344
rect 2684 3336 2692 3344
rect 2636 3276 2644 3284
rect 2604 3176 2612 3184
rect 2588 3076 2596 3084
rect 2588 3056 2596 3064
rect 2668 3216 2676 3224
rect 2636 3136 2644 3144
rect 2636 3096 2644 3104
rect 2668 3096 2676 3104
rect 2668 3076 2676 3084
rect 2668 2896 2676 2904
rect 2588 2836 2596 2844
rect 2668 2756 2676 2764
rect 2652 2716 2660 2724
rect 2540 2676 2548 2684
rect 2572 2676 2580 2684
rect 2508 2596 2516 2604
rect 2492 2576 2500 2584
rect 2444 2496 2452 2504
rect 2476 2496 2484 2504
rect 2316 2296 2324 2304
rect 2444 2296 2452 2304
rect 2348 2276 2356 2284
rect 2396 2276 2404 2284
rect 2380 2256 2388 2264
rect 2428 2256 2436 2264
rect 2204 2116 2212 2124
rect 2188 2096 2196 2104
rect 2252 2136 2260 2144
rect 2316 2156 2324 2164
rect 2268 2116 2276 2124
rect 2300 2116 2308 2124
rect 2252 2096 2260 2104
rect 2172 2056 2180 2064
rect 2236 2056 2244 2064
rect 2124 1936 2132 1944
rect 1980 1916 1988 1924
rect 2012 1916 2020 1924
rect 1868 1876 1876 1884
rect 1900 1876 1908 1884
rect 1916 1876 1924 1884
rect 1788 1816 1796 1824
rect 1852 1816 1860 1824
rect 1836 1796 1844 1804
rect 1788 1716 1796 1724
rect 1884 1716 1892 1724
rect 1820 1676 1828 1684
rect 1868 1676 1876 1684
rect 1676 1656 1684 1664
rect 1708 1656 1716 1664
rect 1756 1656 1764 1664
rect 1660 1636 1668 1644
rect 1708 1636 1716 1644
rect 1564 1576 1572 1584
rect 1564 1496 1572 1504
rect 1596 1496 1604 1504
rect 1500 1476 1508 1484
rect 1484 1456 1492 1464
rect 1404 1356 1412 1364
rect 1388 1236 1396 1244
rect 1548 1476 1556 1484
rect 1532 1456 1540 1464
rect 1516 1436 1524 1444
rect 1612 1456 1620 1464
rect 1580 1396 1588 1404
rect 1596 1396 1604 1404
rect 1916 1676 1924 1684
rect 1900 1616 1908 1624
rect 2124 1916 2132 1924
rect 2076 1896 2084 1904
rect 2188 2016 2196 2024
rect 2156 1896 2164 1904
rect 2236 1896 2244 1904
rect 2252 1896 2260 1904
rect 2284 1896 2292 1904
rect 1980 1876 1988 1884
rect 1964 1856 1972 1864
rect 1980 1856 1988 1864
rect 1948 1836 1956 1844
rect 2060 1836 2068 1844
rect 2076 1836 2084 1844
rect 1964 1796 1972 1804
rect 1996 1756 2004 1764
rect 1964 1716 1972 1724
rect 1996 1716 2004 1724
rect 1932 1636 1940 1644
rect 2172 1856 2180 1864
rect 2092 1816 2100 1824
rect 2108 1816 2116 1824
rect 2236 1816 2244 1824
rect 2268 1876 2276 1884
rect 2284 1776 2292 1784
rect 2252 1736 2260 1744
rect 2108 1716 2116 1724
rect 2060 1696 2068 1704
rect 2044 1676 2052 1684
rect 2124 1656 2132 1664
rect 1996 1636 2004 1644
rect 1788 1516 1796 1524
rect 1836 1516 1844 1524
rect 1724 1496 1732 1504
rect 1804 1496 1812 1504
rect 1868 1496 1876 1504
rect 1932 1496 1940 1504
rect 1948 1496 1956 1504
rect 1740 1476 1748 1484
rect 1868 1476 1876 1484
rect 1900 1476 1908 1484
rect 1756 1436 1764 1444
rect 1660 1376 1668 1384
rect 1596 1356 1604 1364
rect 1612 1356 1620 1364
rect 1388 1216 1396 1224
rect 1484 1216 1492 1224
rect 1411 1206 1419 1214
rect 1421 1206 1429 1214
rect 1431 1206 1439 1214
rect 1441 1206 1449 1214
rect 1451 1206 1459 1214
rect 1461 1206 1469 1214
rect 1308 1196 1316 1204
rect 1356 1196 1364 1204
rect 1388 1196 1396 1204
rect 1260 1096 1268 1104
rect 1276 1076 1284 1084
rect 1244 1056 1252 1064
rect 1292 1036 1300 1044
rect 1276 976 1284 984
rect 1372 1076 1380 1084
rect 1340 1016 1348 1024
rect 1932 1456 1940 1464
rect 1884 1356 1892 1364
rect 1804 1336 1812 1344
rect 1820 1336 1828 1344
rect 1756 1316 1764 1324
rect 1612 1296 1620 1304
rect 1628 1296 1636 1304
rect 1612 1216 1620 1224
rect 1596 1196 1604 1204
rect 1532 1156 1540 1164
rect 1436 1096 1444 1104
rect 1404 1056 1412 1064
rect 1516 1076 1524 1084
rect 1564 1096 1572 1104
rect 1644 1216 1652 1224
rect 1740 1116 1748 1124
rect 1772 1116 1780 1124
rect 1660 1096 1668 1104
rect 1724 1076 1732 1084
rect 1868 1296 1876 1304
rect 1884 1296 1892 1304
rect 1900 1216 1908 1224
rect 1884 1116 1892 1124
rect 1836 1076 1844 1084
rect 1516 1056 1524 1064
rect 1772 1056 1780 1064
rect 1788 1056 1796 1064
rect 1420 1036 1428 1044
rect 1516 1036 1524 1044
rect 1228 956 1236 964
rect 1308 956 1316 964
rect 1276 936 1284 944
rect 1180 916 1188 924
rect 1260 916 1268 924
rect 1612 1036 1620 1044
rect 1660 1036 1668 1044
rect 1532 1016 1540 1024
rect 1852 1056 1860 1064
rect 1676 1016 1684 1024
rect 1820 1016 1828 1024
rect 1836 996 1844 1004
rect 1740 956 1748 964
rect 1932 1336 1940 1344
rect 1948 1196 1956 1204
rect 1916 1076 1924 1084
rect 1948 1056 1956 1064
rect 1932 1016 1940 1024
rect 1900 996 1908 1004
rect 1276 836 1284 844
rect 1164 776 1172 784
rect 1132 756 1140 764
rect 1180 716 1188 724
rect 1324 796 1332 804
rect 1436 916 1444 924
rect 1548 916 1556 924
rect 1388 876 1396 884
rect 1411 806 1419 814
rect 1421 806 1429 814
rect 1431 806 1439 814
rect 1441 806 1449 814
rect 1451 806 1459 814
rect 1461 806 1469 814
rect 1340 756 1348 764
rect 1516 756 1524 764
rect 1340 736 1348 744
rect 1292 716 1300 724
rect 1324 716 1332 724
rect 1228 696 1236 704
rect 1244 696 1252 704
rect 1116 676 1124 684
rect 1148 656 1156 664
rect 1084 576 1092 584
rect 1292 616 1300 624
rect 1260 556 1268 564
rect 940 376 948 384
rect 1084 376 1092 384
rect 924 356 932 364
rect 860 276 868 284
rect 812 216 820 224
rect 908 276 916 284
rect 924 216 932 224
rect 764 176 772 184
rect 876 176 884 184
rect 908 176 916 184
rect 604 156 612 164
rect 684 156 692 164
rect 732 156 740 164
rect 796 156 804 164
rect 572 136 580 144
rect 988 356 996 364
rect 956 336 964 344
rect 956 316 964 324
rect 1116 336 1124 344
rect 1004 316 1012 324
rect 1020 296 1028 304
rect 1148 316 1156 324
rect 1132 256 1140 264
rect 972 236 980 244
rect 1020 236 1028 244
rect 1180 316 1188 324
rect 1180 296 1188 304
rect 1292 536 1300 544
rect 1308 536 1316 544
rect 1228 516 1236 524
rect 1276 516 1284 524
rect 1532 716 1540 724
rect 1356 696 1364 704
rect 1500 696 1508 704
rect 1468 676 1476 684
rect 1340 656 1348 664
rect 1356 616 1364 624
rect 1356 596 1364 604
rect 1388 576 1396 584
rect 1628 736 1636 744
rect 1660 736 1668 744
rect 1612 716 1620 724
rect 1628 716 1636 724
rect 1548 676 1556 684
rect 1596 676 1604 684
rect 1628 676 1636 684
rect 1692 696 1700 704
rect 1580 656 1588 664
rect 1628 656 1636 664
rect 1516 596 1524 604
rect 1628 596 1636 604
rect 1660 596 1668 604
rect 1484 556 1492 564
rect 1532 556 1540 564
rect 1644 536 1652 544
rect 1276 476 1284 484
rect 1260 336 1268 344
rect 1404 516 1412 524
rect 1356 496 1364 504
rect 1340 476 1348 484
rect 1500 476 1508 484
rect 1468 456 1476 464
rect 1411 406 1419 414
rect 1421 406 1429 414
rect 1431 406 1439 414
rect 1441 406 1449 414
rect 1451 406 1459 414
rect 1461 406 1469 414
rect 1340 356 1348 364
rect 1388 356 1396 364
rect 1404 316 1412 324
rect 1212 296 1220 304
rect 1260 296 1268 304
rect 1340 296 1348 304
rect 1228 276 1236 284
rect 1212 256 1220 264
rect 1228 256 1236 264
rect 1164 236 1172 244
rect 1084 196 1092 204
rect 1004 176 1012 184
rect 1020 156 1028 164
rect 1228 156 1236 164
rect 1292 236 1300 244
rect 1324 196 1332 204
rect 1420 276 1428 284
rect 1436 216 1444 224
rect 1308 176 1316 184
rect 1756 916 1764 924
rect 1820 876 1828 884
rect 1868 876 1876 884
rect 1900 876 1908 884
rect 1788 776 1796 784
rect 2012 1616 2020 1624
rect 2220 1716 2228 1724
rect 2268 1716 2276 1724
rect 2188 1696 2196 1704
rect 2220 1696 2228 1704
rect 2172 1676 2180 1684
rect 2156 1516 2164 1524
rect 2044 1496 2052 1504
rect 2012 1396 2020 1404
rect 1996 1316 2004 1324
rect 1980 1196 1988 1204
rect 2028 1356 2036 1364
rect 2028 1296 2036 1304
rect 2044 1296 2052 1304
rect 2092 1476 2100 1484
rect 2076 1456 2084 1464
rect 2076 1356 2084 1364
rect 2156 1396 2164 1404
rect 2124 1340 2132 1344
rect 2124 1336 2132 1340
rect 2140 1336 2148 1344
rect 2140 1316 2148 1324
rect 2252 1496 2260 1504
rect 2236 1456 2244 1464
rect 2204 1376 2212 1384
rect 2188 1356 2196 1364
rect 2188 1336 2196 1344
rect 2060 1256 2068 1264
rect 2060 1216 2068 1224
rect 1996 1016 2004 1024
rect 2028 996 2036 1004
rect 1980 936 1988 944
rect 2092 1076 2100 1084
rect 2076 1056 2084 1064
rect 2124 1056 2132 1064
rect 2076 996 2084 1004
rect 2220 1316 2228 1324
rect 2172 1296 2180 1304
rect 2188 1196 2196 1204
rect 2252 1356 2260 1364
rect 2236 1176 2244 1184
rect 2236 1156 2244 1164
rect 2204 1116 2212 1124
rect 2156 976 2164 984
rect 2060 856 2068 864
rect 2108 876 2116 884
rect 2140 876 2148 884
rect 1996 816 2004 824
rect 2092 816 2100 824
rect 1964 776 1972 784
rect 1948 736 1956 744
rect 1772 716 1780 724
rect 1948 716 1956 724
rect 1980 716 1988 724
rect 1948 696 1956 704
rect 1852 676 1860 684
rect 1708 636 1716 644
rect 2156 856 2164 864
rect 2188 1016 2196 1024
rect 2204 996 2212 1004
rect 2188 976 2196 984
rect 2252 976 2260 984
rect 2332 2140 2340 2144
rect 2332 2136 2340 2140
rect 2332 1996 2340 2004
rect 2316 1896 2324 1904
rect 2492 2356 2500 2364
rect 2508 2336 2516 2344
rect 2540 2636 2548 2644
rect 2732 3196 2740 3204
rect 2844 3556 2852 3564
rect 2860 3536 2868 3544
rect 3036 4116 3044 4124
rect 3036 4076 3044 4084
rect 3292 4836 3300 4844
rect 3420 5236 3428 5244
rect 3484 5296 3492 5304
rect 3564 5296 3572 5304
rect 3436 5156 3444 5164
rect 3436 5136 3444 5144
rect 3356 5116 3364 5124
rect 3372 5102 3380 5104
rect 3372 5096 3380 5102
rect 3468 5236 3476 5244
rect 3452 5076 3460 5084
rect 3436 5056 3444 5064
rect 3484 5116 3492 5124
rect 3484 5096 3492 5104
rect 3564 5096 3572 5104
rect 3532 5076 3540 5084
rect 3356 5016 3364 5024
rect 3388 4996 3396 5004
rect 3404 4916 3412 4924
rect 3340 4856 3348 4864
rect 3388 4856 3396 4864
rect 3308 4736 3316 4744
rect 3388 4696 3396 4704
rect 3516 5036 3524 5044
rect 3468 4936 3476 4944
rect 3548 5016 3556 5024
rect 3612 5416 3620 5424
rect 3644 5416 3652 5424
rect 3724 5376 3732 5384
rect 3596 5296 3604 5304
rect 3596 5116 3604 5124
rect 3580 4976 3588 4984
rect 3532 4936 3540 4944
rect 3532 4916 3540 4924
rect 3580 4916 3588 4924
rect 3468 4896 3476 4904
rect 3452 4836 3460 4844
rect 3452 4796 3460 4804
rect 3484 4876 3492 4884
rect 3612 5036 3620 5044
rect 5923 5406 5931 5414
rect 5933 5406 5941 5414
rect 5943 5406 5951 5414
rect 5953 5406 5961 5414
rect 5963 5406 5971 5414
rect 5973 5406 5981 5414
rect 4316 5396 4324 5404
rect 6924 5396 6932 5404
rect 7052 5396 7060 5404
rect 3916 5376 3924 5384
rect 4396 5376 4404 5384
rect 4556 5376 4564 5384
rect 5436 5376 5444 5384
rect 5628 5376 5636 5384
rect 5756 5376 5764 5384
rect 5852 5376 5860 5384
rect 6492 5376 6500 5384
rect 6604 5376 6612 5384
rect 6796 5376 6804 5384
rect 4204 5356 4212 5364
rect 4316 5356 4324 5364
rect 3852 5336 3860 5344
rect 3948 5336 3956 5344
rect 3948 5296 3956 5304
rect 3996 5296 4004 5304
rect 4012 5116 4020 5124
rect 3740 5102 3748 5104
rect 3740 5096 3748 5102
rect 3964 5096 3972 5104
rect 3676 4956 3684 4964
rect 3676 4936 3684 4944
rect 3596 4896 3604 4904
rect 3628 4896 3636 4904
rect 3564 4796 3572 4804
rect 3420 4776 3428 4784
rect 3436 4776 3444 4784
rect 3564 4756 3572 4764
rect 3404 4676 3412 4684
rect 3388 4656 3396 4664
rect 3212 4636 3220 4644
rect 3308 4636 3316 4644
rect 3228 4596 3236 4604
rect 3164 4576 3172 4584
rect 3292 4536 3300 4544
rect 3180 4436 3188 4444
rect 3196 4436 3204 4444
rect 3228 4436 3236 4444
rect 3100 4416 3108 4424
rect 3148 4416 3156 4424
rect 3084 4356 3092 4364
rect 3180 4256 3188 4264
rect 3100 4216 3108 4224
rect 3084 4096 3092 4104
rect 3148 4096 3156 4104
rect 3068 4076 3076 4084
rect 3052 4056 3060 4064
rect 3036 3996 3044 4004
rect 3084 3956 3092 3964
rect 3036 3916 3044 3924
rect 3036 3896 3044 3904
rect 3132 3896 3140 3904
rect 3260 4316 3268 4324
rect 3292 4316 3300 4324
rect 3228 4216 3236 4224
rect 3404 4596 3412 4604
rect 3356 4536 3364 4544
rect 3356 4496 3364 4504
rect 3324 4436 3332 4444
rect 3564 4676 3572 4684
rect 3500 4636 3508 4644
rect 3452 4616 3460 4624
rect 3484 4596 3492 4604
rect 3468 4556 3476 4564
rect 3532 4596 3540 4604
rect 3660 4916 3668 4924
rect 3692 4876 3700 4884
rect 3708 4776 3716 4784
rect 3580 4616 3588 4624
rect 3644 4616 3652 4624
rect 3580 4596 3588 4604
rect 3548 4576 3556 4584
rect 3564 4576 3572 4584
rect 3500 4556 3508 4564
rect 3532 4556 3540 4564
rect 3548 4556 3556 4564
rect 3484 4536 3492 4544
rect 3484 4516 3492 4524
rect 3452 4496 3460 4504
rect 3420 4396 3428 4404
rect 3436 4396 3444 4404
rect 3324 4316 3332 4324
rect 3388 4296 3396 4304
rect 3452 4316 3460 4324
rect 3820 4916 3828 4924
rect 3804 4796 3812 4804
rect 3980 5076 3988 5084
rect 4108 5316 4116 5324
rect 4652 5336 4660 5344
rect 4252 5316 4260 5324
rect 4348 5316 4356 5324
rect 4508 5316 4516 5324
rect 4588 5316 4596 5324
rect 4236 5256 4244 5264
rect 4300 5256 4308 5264
rect 4204 5236 4212 5244
rect 4108 5096 4116 5104
rect 3852 4836 3860 4844
rect 4044 5036 4052 5044
rect 4012 4996 4020 5004
rect 3916 4936 3924 4944
rect 3964 4936 3972 4944
rect 3900 4896 3908 4904
rect 3948 4856 3956 4864
rect 3932 4836 3940 4844
rect 3868 4816 3876 4824
rect 3692 4656 3700 4664
rect 3836 4656 3844 4664
rect 3676 4576 3684 4584
rect 3612 4556 3620 4564
rect 3644 4556 3652 4564
rect 3564 4516 3572 4524
rect 3596 4496 3604 4504
rect 3708 4616 3716 4624
rect 3772 4576 3780 4584
rect 3692 4556 3700 4564
rect 3644 4536 3652 4544
rect 3628 4336 3636 4344
rect 3532 4316 3540 4324
rect 3436 4296 3444 4304
rect 3340 4276 3348 4284
rect 3404 4276 3412 4284
rect 3420 4276 3428 4284
rect 3292 4136 3300 4144
rect 3388 4136 3396 4144
rect 3468 4156 3476 4164
rect 3468 4136 3476 4144
rect 3244 4116 3252 4124
rect 3228 4096 3236 4104
rect 3212 3976 3220 3984
rect 3196 3956 3204 3964
rect 3212 3956 3220 3964
rect 3180 3896 3188 3904
rect 3052 3876 3060 3884
rect 3164 3856 3172 3864
rect 3148 3836 3156 3844
rect 3052 3776 3060 3784
rect 3036 3736 3044 3744
rect 3036 3696 3044 3704
rect 2844 3476 2852 3484
rect 3020 3476 3028 3484
rect 2860 3376 2868 3384
rect 2780 3196 2788 3204
rect 2828 3196 2836 3204
rect 2828 3156 2836 3164
rect 2764 3116 2772 3124
rect 2828 3096 2836 3104
rect 2796 3076 2804 3084
rect 2780 3036 2788 3044
rect 2748 2996 2756 3004
rect 2748 2956 2756 2964
rect 2812 2976 2820 2984
rect 2700 2896 2708 2904
rect 2876 3016 2884 3024
rect 2876 2976 2884 2984
rect 2915 3406 2923 3414
rect 2925 3406 2933 3414
rect 2935 3406 2943 3414
rect 2945 3406 2953 3414
rect 2955 3406 2963 3414
rect 2965 3406 2973 3414
rect 2972 3376 2980 3384
rect 2940 3356 2948 3364
rect 3324 4036 3332 4044
rect 3260 3856 3268 3864
rect 3292 3856 3300 3864
rect 3228 3836 3236 3844
rect 3260 3836 3268 3844
rect 3100 3776 3108 3784
rect 3212 3776 3220 3784
rect 3228 3736 3236 3744
rect 3068 3676 3076 3684
rect 3180 3676 3188 3684
rect 3100 3516 3108 3524
rect 3068 3436 3076 3444
rect 3148 3476 3156 3484
rect 3244 3476 3252 3484
rect 3132 3416 3140 3424
rect 3324 3876 3332 3884
rect 3324 3856 3332 3864
rect 3308 3716 3316 3724
rect 3356 3756 3364 3764
rect 3340 3736 3348 3744
rect 3356 3716 3364 3724
rect 3436 4076 3444 4084
rect 3532 4236 3540 4244
rect 3516 4216 3524 4224
rect 3500 4136 3508 4144
rect 3484 4116 3492 4124
rect 3452 3996 3460 4004
rect 3436 3976 3444 3984
rect 3468 3976 3476 3984
rect 3468 3956 3476 3964
rect 3436 3876 3444 3884
rect 3388 3776 3396 3784
rect 3340 3696 3348 3704
rect 3324 3656 3332 3664
rect 3404 3716 3412 3724
rect 3452 3716 3460 3724
rect 3420 3696 3428 3704
rect 3436 3676 3444 3684
rect 3452 3676 3460 3684
rect 3500 4096 3508 4104
rect 3548 4136 3556 4144
rect 3564 4056 3572 4064
rect 3532 3976 3540 3984
rect 3564 3836 3572 3844
rect 3500 3776 3508 3784
rect 3516 3776 3524 3784
rect 3500 3736 3508 3744
rect 3516 3676 3524 3684
rect 3484 3616 3492 3624
rect 3548 3696 3556 3704
rect 3436 3596 3444 3604
rect 3532 3596 3540 3604
rect 3292 3516 3300 3524
rect 3276 3416 3284 3424
rect 3196 3356 3204 3364
rect 2908 3296 2916 3304
rect 3084 3276 3092 3284
rect 3052 3256 3060 3264
rect 3116 3256 3124 3264
rect 3100 3236 3108 3244
rect 3020 3176 3028 3184
rect 3004 3156 3012 3164
rect 2988 3116 2996 3124
rect 2972 3056 2980 3064
rect 2915 3006 2923 3014
rect 2925 3006 2933 3014
rect 2935 3006 2943 3014
rect 2945 3006 2953 3014
rect 2955 3006 2963 3014
rect 2965 3006 2973 3014
rect 2892 2956 2900 2964
rect 2892 2936 2900 2944
rect 2940 2936 2948 2944
rect 2908 2916 2916 2924
rect 2844 2896 2852 2904
rect 2828 2876 2836 2884
rect 2876 2876 2884 2884
rect 2780 2796 2788 2804
rect 2700 2716 2708 2724
rect 2684 2696 2692 2704
rect 2716 2696 2724 2704
rect 2652 2676 2660 2684
rect 2716 2676 2724 2684
rect 2860 2736 2868 2744
rect 3052 3156 3060 3164
rect 3052 3136 3060 3144
rect 3036 3056 3044 3064
rect 3292 3356 3300 3364
rect 3212 3216 3220 3224
rect 3356 3476 3364 3484
rect 3484 3576 3492 3584
rect 3452 3516 3460 3524
rect 3372 3456 3380 3464
rect 3388 3456 3396 3464
rect 3404 3456 3412 3464
rect 3420 3456 3428 3464
rect 3596 4276 3604 4284
rect 3756 4516 3764 4524
rect 3756 4496 3764 4504
rect 3692 4336 3700 4344
rect 3644 4316 3652 4324
rect 3724 4456 3732 4464
rect 3804 4516 3812 4524
rect 3836 4476 3844 4484
rect 3884 4556 3892 4564
rect 3868 4456 3876 4464
rect 3788 4396 3796 4404
rect 3708 4296 3716 4304
rect 3628 4196 3636 4204
rect 3612 4136 3620 4144
rect 3724 4276 3732 4284
rect 3708 4256 3716 4264
rect 3740 4216 3748 4224
rect 3740 4176 3748 4184
rect 3692 4136 3700 4144
rect 3708 4136 3716 4144
rect 3612 4116 3620 4124
rect 3676 4116 3684 4124
rect 3740 4116 3748 4124
rect 3676 4016 3684 4024
rect 3788 4176 3796 4184
rect 3756 4036 3764 4044
rect 3724 3956 3732 3964
rect 3596 3902 3604 3904
rect 3596 3896 3604 3902
rect 3660 3896 3668 3904
rect 3580 3796 3588 3804
rect 3900 4516 3908 4524
rect 3932 4476 3940 4484
rect 3916 4456 3924 4464
rect 4419 5206 4427 5214
rect 4429 5206 4437 5214
rect 4439 5206 4447 5214
rect 4449 5206 4457 5214
rect 4459 5206 4467 5214
rect 4469 5206 4477 5214
rect 4236 5116 4244 5124
rect 4380 5116 4388 5124
rect 4268 5096 4276 5104
rect 4204 5036 4212 5044
rect 4220 5036 4228 5044
rect 4140 4956 4148 4964
rect 4060 4936 4068 4944
rect 4284 5076 4292 5084
rect 4252 5056 4260 5064
rect 4332 5096 4340 5104
rect 4364 5076 4372 5084
rect 4460 5076 4468 5084
rect 4300 5056 4308 5064
rect 4332 5036 4340 5044
rect 4428 5036 4436 5044
rect 4252 4976 4260 4984
rect 4444 4976 4452 4984
rect 4236 4936 4244 4944
rect 4188 4856 4196 4864
rect 3996 4836 4004 4844
rect 4076 4836 4084 4844
rect 4108 4716 4116 4724
rect 4236 4716 4244 4724
rect 3996 4702 4004 4704
rect 3996 4696 4004 4702
rect 4076 4676 4084 4684
rect 3964 4576 3972 4584
rect 4028 4556 4036 4564
rect 3980 4516 3988 4524
rect 4012 4516 4020 4524
rect 4092 4556 4100 4564
rect 4332 4936 4340 4944
rect 4348 4936 4356 4944
rect 4396 4936 4404 4944
rect 4316 4836 4324 4844
rect 4124 4696 4132 4704
rect 4204 4696 4212 4704
rect 4284 4696 4292 4704
rect 4300 4696 4308 4704
rect 4156 4676 4164 4684
rect 4364 4736 4372 4744
rect 4348 4696 4356 4704
rect 4332 4676 4340 4684
rect 4188 4656 4196 4664
rect 4236 4656 4244 4664
rect 4172 4636 4180 4644
rect 4284 4576 4292 4584
rect 4156 4556 4164 4564
rect 4108 4536 4116 4544
rect 4188 4536 4196 4544
rect 4236 4536 4244 4544
rect 4060 4496 4068 4504
rect 3964 4476 3972 4484
rect 3948 4416 3956 4424
rect 3948 4396 3956 4404
rect 3996 4456 4004 4464
rect 4012 4376 4020 4384
rect 4316 4656 4324 4664
rect 4492 4856 4500 4864
rect 4419 4806 4427 4814
rect 4429 4806 4437 4814
rect 4439 4806 4447 4814
rect 4449 4806 4457 4814
rect 4459 4806 4467 4814
rect 4469 4806 4477 4814
rect 4540 5176 4548 5184
rect 5292 5356 5300 5364
rect 5340 5356 5348 5364
rect 5564 5356 5572 5364
rect 4796 5336 4804 5344
rect 5260 5336 5268 5344
rect 4700 5316 4708 5324
rect 4620 5256 4628 5264
rect 4668 5256 4676 5264
rect 4636 5216 4644 5224
rect 4572 5156 4580 5164
rect 4556 5056 4564 5064
rect 4620 5116 4628 5124
rect 4604 5076 4612 5084
rect 4588 5036 4596 5044
rect 4620 5036 4628 5044
rect 4572 4996 4580 5004
rect 4556 4956 4564 4964
rect 4572 4956 4580 4964
rect 4540 4896 4548 4904
rect 4604 4996 4612 5004
rect 4604 4896 4612 4904
rect 4588 4856 4596 4864
rect 4524 4816 4532 4824
rect 4508 4776 4516 4784
rect 4524 4736 4532 4744
rect 4492 4716 4500 4724
rect 4508 4696 4516 4704
rect 4332 4556 4340 4564
rect 4396 4556 4404 4564
rect 4268 4516 4276 4524
rect 4300 4516 4308 4524
rect 4476 4516 4484 4524
rect 4028 4356 4036 4364
rect 4156 4302 4164 4304
rect 4156 4296 4164 4302
rect 4188 4296 4196 4304
rect 3964 4256 3972 4264
rect 4156 4256 4164 4264
rect 3820 4176 3828 4184
rect 3980 4176 3988 4184
rect 3884 4136 3892 4144
rect 3948 4136 3956 4144
rect 3868 4116 3876 4124
rect 3820 4076 3828 4084
rect 4092 4216 4100 4224
rect 4236 4276 4244 4284
rect 4028 4196 4036 4204
rect 4076 4176 4084 4184
rect 4108 4156 4116 4164
rect 4188 4156 4196 4164
rect 4012 4076 4020 4084
rect 4012 4036 4020 4044
rect 3820 3976 3828 3984
rect 3916 3916 3924 3924
rect 3804 3876 3812 3884
rect 3868 3876 3876 3884
rect 3740 3856 3748 3864
rect 3596 3776 3604 3784
rect 3724 3776 3732 3784
rect 3788 3836 3796 3844
rect 3852 3796 3860 3804
rect 3772 3776 3780 3784
rect 3836 3776 3844 3784
rect 3676 3756 3684 3764
rect 3756 3756 3764 3764
rect 3580 3676 3588 3684
rect 3708 3736 3716 3744
rect 3804 3756 3812 3764
rect 3820 3756 3828 3764
rect 3852 3756 3860 3764
rect 3692 3716 3700 3724
rect 3740 3716 3748 3724
rect 3820 3716 3828 3724
rect 3756 3696 3764 3704
rect 3740 3656 3748 3664
rect 3612 3636 3620 3644
rect 3596 3516 3604 3524
rect 3468 3496 3476 3504
rect 3468 3476 3476 3484
rect 3516 3476 3524 3484
rect 3596 3476 3604 3484
rect 3452 3436 3460 3444
rect 3388 3376 3396 3384
rect 3340 3356 3348 3364
rect 3324 3316 3332 3324
rect 3452 3316 3460 3324
rect 3484 3456 3492 3464
rect 3500 3416 3508 3424
rect 3484 3296 3492 3304
rect 3404 3276 3412 3284
rect 3308 3196 3316 3204
rect 3132 2976 3140 2984
rect 3068 2956 3076 2964
rect 3292 3036 3300 3044
rect 3212 2996 3220 3004
rect 3276 2956 3284 2964
rect 3228 2936 3236 2944
rect 3196 2916 3204 2924
rect 3340 3136 3348 3144
rect 3308 2916 3316 2924
rect 3084 2896 3092 2904
rect 3148 2896 3156 2904
rect 3212 2896 3220 2904
rect 3180 2876 3188 2884
rect 3244 2876 3252 2884
rect 3388 3256 3396 3264
rect 3436 3256 3444 3264
rect 3452 3256 3460 3264
rect 3420 3216 3428 3224
rect 3452 3156 3460 3164
rect 3404 3096 3412 3104
rect 3548 3456 3556 3464
rect 3724 3556 3732 3564
rect 3756 3576 3764 3584
rect 3788 3516 3796 3524
rect 3788 3496 3796 3504
rect 3676 3476 3684 3484
rect 3708 3480 3716 3484
rect 3708 3476 3716 3480
rect 3740 3456 3748 3464
rect 3820 3556 3828 3564
rect 3932 3856 3940 3864
rect 3884 3836 3892 3844
rect 3900 3796 3908 3804
rect 3996 3736 4004 3744
rect 3852 3716 3860 3724
rect 3868 3716 3876 3724
rect 3868 3616 3876 3624
rect 3836 3496 3844 3504
rect 3644 3436 3652 3444
rect 3740 3436 3748 3444
rect 3676 3396 3684 3404
rect 3532 3356 3540 3364
rect 3548 3356 3556 3364
rect 3644 3356 3652 3364
rect 3708 3356 3716 3364
rect 3516 3336 3524 3344
rect 3564 3336 3572 3344
rect 3580 3316 3588 3324
rect 3612 3316 3620 3324
rect 3708 3316 3716 3324
rect 3772 3318 3780 3324
rect 3772 3316 3780 3318
rect 3660 3296 3668 3304
rect 3548 3276 3556 3284
rect 3724 3276 3732 3284
rect 3612 3256 3620 3264
rect 3628 3196 3636 3204
rect 3468 3136 3476 3144
rect 3532 3136 3540 3144
rect 3644 3136 3652 3144
rect 3708 3136 3716 3144
rect 3468 3096 3476 3104
rect 3516 3096 3524 3104
rect 3404 3076 3412 3084
rect 3436 3056 3444 3064
rect 3420 2976 3428 2984
rect 3388 2956 3396 2964
rect 3356 2936 3364 2944
rect 3340 2896 3348 2904
rect 3260 2856 3268 2864
rect 3052 2816 3060 2824
rect 2780 2696 2788 2704
rect 2860 2696 2868 2704
rect 2764 2676 2772 2684
rect 2732 2656 2740 2664
rect 2828 2656 2836 2664
rect 2492 2236 2500 2244
rect 2540 2316 2548 2324
rect 2572 2376 2580 2384
rect 2668 2316 2676 2324
rect 2556 2276 2564 2284
rect 2716 2516 2724 2524
rect 2700 2436 2708 2444
rect 2540 2256 2548 2264
rect 2524 2216 2532 2224
rect 2604 2216 2612 2224
rect 2620 2216 2628 2224
rect 2620 2176 2628 2184
rect 2636 2176 2644 2184
rect 2684 2256 2692 2264
rect 2700 2256 2708 2264
rect 2684 2176 2692 2184
rect 2764 2476 2772 2484
rect 2748 2356 2756 2364
rect 2748 2296 2756 2304
rect 2748 2276 2756 2284
rect 2748 2176 2756 2184
rect 2460 2156 2468 2164
rect 2540 2156 2548 2164
rect 2668 2156 2676 2164
rect 2748 2156 2756 2164
rect 2460 2136 2468 2144
rect 2364 2116 2372 2124
rect 2428 2096 2436 2104
rect 2364 2056 2372 2064
rect 2412 2056 2420 2064
rect 2380 2036 2388 2044
rect 2396 2036 2404 2044
rect 2348 1956 2356 1964
rect 2364 1916 2372 1924
rect 2396 1936 2404 1944
rect 2444 2056 2452 2064
rect 2428 1856 2436 1864
rect 2396 1836 2404 1844
rect 2412 1776 2420 1784
rect 2348 1736 2356 1744
rect 2396 1716 2404 1724
rect 2348 1656 2356 1664
rect 2396 1696 2404 1704
rect 2364 1636 2372 1644
rect 2460 2016 2468 2024
rect 2508 2016 2516 2024
rect 2572 2136 2580 2144
rect 2668 2116 2676 2124
rect 2716 2116 2724 2124
rect 2556 2096 2564 2104
rect 2636 2096 2644 2104
rect 2732 2096 2740 2104
rect 2540 1936 2548 1944
rect 2492 1916 2500 1924
rect 2524 1836 2532 1844
rect 2604 1916 2612 1924
rect 2556 1876 2564 1884
rect 2460 1776 2468 1784
rect 2492 1756 2500 1764
rect 2460 1696 2468 1704
rect 2508 1676 2516 1684
rect 2540 1696 2548 1704
rect 2524 1656 2532 1664
rect 2604 1836 2612 1844
rect 2620 1836 2628 1844
rect 2572 1736 2580 1744
rect 2620 1736 2628 1744
rect 2604 1716 2612 1724
rect 2572 1696 2580 1704
rect 2620 1536 2628 1544
rect 2348 1516 2356 1524
rect 2444 1516 2452 1524
rect 2316 1456 2324 1464
rect 2284 1436 2292 1444
rect 2332 1436 2340 1444
rect 2412 1496 2420 1504
rect 2476 1496 2484 1504
rect 2572 1496 2580 1504
rect 2364 1476 2372 1484
rect 2364 1456 2372 1464
rect 2364 1376 2372 1384
rect 2284 1336 2292 1344
rect 2348 1356 2356 1364
rect 2428 1476 2436 1484
rect 2428 1456 2436 1464
rect 2444 1456 2452 1464
rect 2556 1456 2564 1464
rect 2524 1436 2532 1444
rect 2460 1396 2468 1404
rect 2492 1396 2500 1404
rect 2380 1316 2388 1324
rect 2332 1296 2340 1304
rect 2364 1256 2372 1264
rect 2396 1256 2404 1264
rect 2444 1256 2452 1264
rect 2348 1096 2356 1104
rect 2300 1076 2308 1084
rect 2332 1056 2340 1064
rect 2284 996 2292 1004
rect 2348 996 2356 1004
rect 2236 916 2244 924
rect 2300 916 2308 924
rect 2268 856 2276 864
rect 2172 816 2180 824
rect 2252 756 2260 764
rect 2316 816 2324 824
rect 2332 816 2340 824
rect 2188 716 2196 724
rect 2236 716 2244 724
rect 1996 696 2004 704
rect 2124 696 2132 704
rect 2188 696 2196 704
rect 2300 736 2308 744
rect 2284 696 2292 704
rect 2156 676 2164 684
rect 2220 676 2228 684
rect 1836 656 1844 664
rect 1740 636 1748 644
rect 1724 596 1732 604
rect 1788 596 1796 604
rect 1836 596 1844 604
rect 1868 596 1876 604
rect 1948 596 1956 604
rect 1724 556 1732 564
rect 1740 556 1748 564
rect 1836 556 1844 564
rect 1708 536 1716 544
rect 1772 536 1780 544
rect 1868 536 1876 544
rect 1596 516 1604 524
rect 1820 516 1828 524
rect 1580 496 1588 504
rect 1548 376 1556 384
rect 1644 476 1652 484
rect 1756 456 1764 464
rect 1612 356 1620 364
rect 1836 336 1844 344
rect 2092 656 2100 664
rect 1996 556 2004 564
rect 2028 556 2036 564
rect 2092 556 2100 564
rect 2140 576 2148 584
rect 2204 616 2212 624
rect 2268 656 2276 664
rect 2156 556 2164 564
rect 2188 556 2196 564
rect 2220 556 2228 564
rect 2252 556 2260 564
rect 2012 536 2020 544
rect 2108 536 2116 544
rect 1916 516 1924 524
rect 1964 516 1972 524
rect 2060 516 2068 524
rect 2156 496 2164 504
rect 1868 376 1876 384
rect 1868 336 1876 344
rect 1596 296 1604 304
rect 1628 316 1636 324
rect 1692 316 1700 324
rect 1852 316 1860 324
rect 1964 376 1972 384
rect 1932 316 1940 324
rect 1708 296 1716 304
rect 1804 296 1812 304
rect 1612 276 1620 284
rect 1596 256 1604 264
rect 1756 256 1764 264
rect 1532 236 1540 244
rect 1516 176 1524 184
rect 1532 176 1540 184
rect 748 136 756 144
rect 860 136 868 144
rect 1116 136 1124 144
rect 1244 136 1252 144
rect 380 116 388 124
rect 444 116 452 124
rect 540 116 548 124
rect 860 116 868 124
rect 908 116 916 124
rect 28 96 36 104
rect 204 96 212 104
rect 284 96 292 104
rect 316 96 324 104
rect 1644 236 1652 244
rect 1612 196 1620 204
rect 1660 216 1668 224
rect 1708 216 1716 224
rect 1660 196 1668 204
rect 1628 156 1636 164
rect 1628 116 1636 124
rect 444 96 452 104
rect 492 96 500 104
rect 604 96 612 104
rect 636 96 644 104
rect 1132 96 1140 104
rect 1548 96 1556 104
rect 1740 156 1748 164
rect 1852 276 1860 284
rect 2028 356 2036 364
rect 1964 256 1972 264
rect 1916 236 1924 244
rect 1884 216 1892 224
rect 1868 196 1876 204
rect 1804 176 1812 184
rect 1692 136 1700 144
rect 1676 116 1684 124
rect 1740 116 1748 124
rect 1820 156 1828 164
rect 1980 236 1988 244
rect 1996 196 2004 204
rect 1996 176 2004 184
rect 2092 316 2100 324
rect 2124 316 2132 324
rect 2140 316 2148 324
rect 2236 516 2244 524
rect 2204 376 2212 384
rect 2236 336 2244 344
rect 2220 316 2228 324
rect 2172 276 2180 284
rect 2188 276 2196 284
rect 2028 256 2036 264
rect 2156 256 2164 264
rect 2092 236 2100 244
rect 2140 236 2148 244
rect 2076 196 2084 204
rect 2108 176 2116 184
rect 2012 156 2020 164
rect 2188 236 2196 244
rect 2300 636 2308 644
rect 2284 596 2292 604
rect 2396 1196 2404 1204
rect 2588 1476 2596 1484
rect 2604 1476 2612 1484
rect 2604 1396 2612 1404
rect 2732 2056 2740 2064
rect 2668 2016 2676 2024
rect 2732 1896 2740 1904
rect 2684 1796 2692 1804
rect 2668 1776 2676 1784
rect 2732 1776 2740 1784
rect 2828 2536 2836 2544
rect 2844 2516 2852 2524
rect 2812 2496 2820 2504
rect 2844 2496 2852 2504
rect 2796 2456 2804 2464
rect 2780 2376 2788 2384
rect 2780 2336 2788 2344
rect 2876 2676 2884 2684
rect 2915 2606 2923 2614
rect 2925 2606 2933 2614
rect 2935 2606 2943 2614
rect 2945 2606 2953 2614
rect 2955 2606 2963 2614
rect 2965 2606 2973 2614
rect 3020 2576 3028 2584
rect 2972 2436 2980 2444
rect 3100 2676 3108 2684
rect 3084 2616 3092 2624
rect 3132 2776 3140 2784
rect 3148 2776 3156 2784
rect 3116 2596 3124 2604
rect 3116 2576 3124 2584
rect 3228 2776 3236 2784
rect 3276 2776 3284 2784
rect 3196 2696 3204 2704
rect 3212 2676 3220 2684
rect 3212 2656 3220 2664
rect 3196 2636 3204 2644
rect 3196 2616 3204 2624
rect 3148 2596 3156 2604
rect 3068 2516 3076 2524
rect 3100 2516 3108 2524
rect 2988 2396 2996 2404
rect 3020 2376 3028 2384
rect 3004 2356 3012 2364
rect 3052 2356 3060 2364
rect 2780 2296 2788 2304
rect 2860 2296 2868 2304
rect 3020 2296 3028 2304
rect 2796 2276 2804 2284
rect 2812 2276 2820 2284
rect 3036 2276 3044 2284
rect 2844 2236 2852 2244
rect 2908 2236 2916 2244
rect 2915 2206 2923 2214
rect 2925 2206 2933 2214
rect 2935 2206 2943 2214
rect 2945 2206 2953 2214
rect 2955 2206 2963 2214
rect 2965 2206 2973 2214
rect 3036 2176 3044 2184
rect 3116 2336 3124 2344
rect 3148 2336 3156 2344
rect 3196 2396 3204 2404
rect 3244 2716 3252 2724
rect 3260 2696 3268 2704
rect 3356 2856 3364 2864
rect 3372 2756 3380 2764
rect 3500 3036 3508 3044
rect 3516 3016 3524 3024
rect 3484 2976 3492 2984
rect 3452 2956 3460 2964
rect 3468 2936 3476 2944
rect 3548 3096 3556 3104
rect 3452 2916 3460 2924
rect 3580 3096 3588 3104
rect 3596 3056 3604 3064
rect 3676 3096 3684 3104
rect 3628 3076 3636 3084
rect 3644 3076 3652 3084
rect 3644 2996 3652 3004
rect 3660 2956 3668 2964
rect 3836 3456 3844 3464
rect 3852 3456 3860 3464
rect 3836 3316 3844 3324
rect 3868 3296 3876 3304
rect 3932 3716 3940 3724
rect 3980 3716 3988 3724
rect 3964 3676 3972 3684
rect 3948 3656 3956 3664
rect 3980 3576 3988 3584
rect 3932 3556 3940 3564
rect 3916 3496 3924 3504
rect 3996 3556 4004 3564
rect 4140 4116 4148 4124
rect 4204 4096 4212 4104
rect 4124 4076 4132 4084
rect 4092 3976 4100 3984
rect 4108 3916 4116 3924
rect 4028 3880 4036 3884
rect 4028 3876 4036 3880
rect 4044 3876 4052 3884
rect 4076 3856 4084 3864
rect 4060 3756 4068 3764
rect 4028 3716 4036 3724
rect 4044 3696 4052 3704
rect 3996 3536 4004 3544
rect 4012 3536 4020 3544
rect 4220 3996 4228 4004
rect 4188 3976 4196 3984
rect 4172 3916 4180 3924
rect 4124 3796 4132 3804
rect 4156 3876 4164 3884
rect 4204 3836 4212 3844
rect 4419 4406 4427 4414
rect 4429 4406 4437 4414
rect 4439 4406 4447 4414
rect 4449 4406 4457 4414
rect 4459 4406 4467 4414
rect 4469 4406 4477 4414
rect 4540 4576 4548 4584
rect 4508 4556 4516 4564
rect 4620 4776 4628 4784
rect 4620 4756 4628 4764
rect 4796 5176 4804 5184
rect 4684 5136 4692 5144
rect 4748 5116 4756 5124
rect 4764 5096 4772 5104
rect 4652 5076 4660 5084
rect 4684 5036 4692 5044
rect 4700 5036 4708 5044
rect 4716 5016 4724 5024
rect 4732 5016 4740 5024
rect 4748 4996 4756 5004
rect 4764 4956 4772 4964
rect 4652 4896 4660 4904
rect 4684 4856 4692 4864
rect 4732 4856 4740 4864
rect 4764 4856 4772 4864
rect 4828 5316 4836 5324
rect 4972 5316 4980 5324
rect 4796 4996 4804 5004
rect 4812 4996 4820 5004
rect 4924 5296 4932 5304
rect 4956 5296 4964 5304
rect 5052 5316 5060 5324
rect 4988 5236 4996 5244
rect 5196 5316 5204 5324
rect 5308 5316 5316 5324
rect 5676 5356 5684 5364
rect 5596 5336 5604 5344
rect 5388 5316 5396 5324
rect 5308 5296 5316 5304
rect 5356 5296 5364 5304
rect 5372 5296 5380 5304
rect 5372 5276 5380 5284
rect 5004 5216 5012 5224
rect 5052 5216 5060 5224
rect 4908 5196 4916 5204
rect 5020 5196 5028 5204
rect 5340 5196 5348 5204
rect 5084 5176 5092 5184
rect 5116 5156 5124 5164
rect 4892 5116 4900 5124
rect 5308 5136 5316 5144
rect 5148 5116 5156 5124
rect 5164 5116 5172 5124
rect 5228 5116 5236 5124
rect 5244 5116 5252 5124
rect 5324 5116 5332 5124
rect 4860 5076 4868 5084
rect 4908 5076 4916 5084
rect 4876 5036 4884 5044
rect 4844 5016 4852 5024
rect 5004 5076 5012 5084
rect 4860 4996 4868 5004
rect 4956 4996 4964 5004
rect 5084 5076 5092 5084
rect 5068 5036 5076 5044
rect 5052 5016 5060 5024
rect 4988 4976 4996 4984
rect 5020 4956 5028 4964
rect 5068 4956 5076 4964
rect 4908 4936 4916 4944
rect 5068 4936 5076 4944
rect 4652 4816 4660 4824
rect 4668 4816 4676 4824
rect 4636 4736 4644 4744
rect 4652 4696 4660 4704
rect 4636 4676 4644 4684
rect 4732 4756 4740 4764
rect 4700 4736 4708 4744
rect 4684 4656 4692 4664
rect 4732 4656 4740 4664
rect 4748 4656 4756 4664
rect 4812 4756 4820 4764
rect 4812 4736 4820 4744
rect 4780 4656 4788 4664
rect 4764 4636 4772 4644
rect 4668 4576 4676 4584
rect 4556 4516 4564 4524
rect 4636 4516 4644 4524
rect 4716 4516 4724 4524
rect 4524 4436 4532 4444
rect 4332 4276 4340 4284
rect 4444 4276 4452 4284
rect 4316 4256 4324 4264
rect 4284 3996 4292 4004
rect 4476 4156 4484 4164
rect 4396 4136 4404 4144
rect 4252 3916 4260 3924
rect 4236 3796 4244 3804
rect 4268 3796 4276 3804
rect 4092 3776 4100 3784
rect 4220 3776 4228 3784
rect 4108 3756 4116 3764
rect 4172 3756 4180 3764
rect 4236 3756 4244 3764
rect 4108 3676 4116 3684
rect 4124 3676 4132 3684
rect 4140 3676 4148 3684
rect 4076 3536 4084 3544
rect 4092 3516 4100 3524
rect 4124 3536 4132 3544
rect 3980 3496 3988 3504
rect 4044 3496 4052 3504
rect 4108 3496 4116 3504
rect 3900 3476 3908 3484
rect 3900 3376 3908 3384
rect 3932 3456 3940 3464
rect 3948 3456 3956 3464
rect 3932 3396 3940 3404
rect 3884 3276 3892 3284
rect 3740 3156 3748 3164
rect 3772 3156 3780 3164
rect 3772 3116 3780 3124
rect 3788 3116 3796 3124
rect 3724 3056 3732 3064
rect 3708 3036 3716 3044
rect 3692 3016 3700 3024
rect 3708 2996 3716 3004
rect 3612 2936 3620 2944
rect 3676 2936 3684 2944
rect 3692 2936 3700 2944
rect 3612 2916 3620 2924
rect 3468 2896 3476 2904
rect 3532 2896 3540 2904
rect 3564 2896 3572 2904
rect 3580 2896 3588 2904
rect 3628 2896 3636 2904
rect 3484 2876 3492 2884
rect 3420 2776 3428 2784
rect 3420 2716 3428 2724
rect 3356 2696 3364 2704
rect 3324 2676 3332 2684
rect 3356 2676 3364 2684
rect 3276 2656 3284 2664
rect 3420 2676 3428 2684
rect 3404 2636 3412 2644
rect 3324 2576 3332 2584
rect 3276 2556 3284 2564
rect 3372 2536 3380 2544
rect 3292 2496 3300 2504
rect 3356 2436 3364 2444
rect 3276 2336 3284 2344
rect 3388 2416 3396 2424
rect 3164 2316 3172 2324
rect 3244 2316 3252 2324
rect 3372 2316 3380 2324
rect 3084 2296 3092 2304
rect 3148 2296 3156 2304
rect 3276 2296 3284 2304
rect 2780 2136 2788 2144
rect 2956 2136 2964 2144
rect 2764 2056 2772 2064
rect 2764 1976 2772 1984
rect 2844 2076 2852 2084
rect 2860 2076 2868 2084
rect 2844 2016 2852 2024
rect 2780 1956 2788 1964
rect 2764 1896 2772 1904
rect 2780 1896 2788 1904
rect 2748 1756 2756 1764
rect 2812 1956 2820 1964
rect 3068 2076 3076 2084
rect 2876 1996 2884 2004
rect 3052 1996 3060 2004
rect 2812 1916 2820 1924
rect 2828 1896 2836 1904
rect 2892 1916 2900 1924
rect 2892 1896 2900 1904
rect 3020 1896 3028 1904
rect 2908 1876 2916 1884
rect 3036 1876 3044 1884
rect 2876 1856 2884 1864
rect 3100 2276 3108 2284
rect 3164 2276 3172 2284
rect 3292 2276 3300 2284
rect 3084 1896 3092 1904
rect 3228 2236 3236 2244
rect 3260 2236 3268 2244
rect 3308 2236 3316 2244
rect 3340 2236 3348 2244
rect 3372 2236 3380 2244
rect 3228 2216 3236 2224
rect 3116 2156 3124 2164
rect 3116 2136 3124 2144
rect 3228 2136 3236 2144
rect 3308 2136 3316 2144
rect 3164 2116 3172 2124
rect 3212 2116 3220 2124
rect 3260 2116 3268 2124
rect 3132 1936 3140 1944
rect 3100 1876 3108 1884
rect 2844 1816 2852 1824
rect 2844 1796 2852 1804
rect 2828 1756 2836 1764
rect 2796 1736 2804 1744
rect 2716 1716 2724 1724
rect 2780 1716 2788 1724
rect 2700 1616 2708 1624
rect 2652 1556 2660 1564
rect 2764 1616 2772 1624
rect 2796 1616 2804 1624
rect 3036 1836 3044 1844
rect 2915 1806 2923 1814
rect 2925 1806 2933 1814
rect 2935 1806 2943 1814
rect 2945 1806 2953 1814
rect 2955 1806 2963 1814
rect 2965 1806 2973 1814
rect 2940 1776 2948 1784
rect 2844 1716 2852 1724
rect 2892 1716 2900 1724
rect 2876 1676 2884 1684
rect 2812 1536 2820 1544
rect 2716 1496 2724 1504
rect 2668 1476 2676 1484
rect 2700 1476 2708 1484
rect 2748 1476 2756 1484
rect 2812 1476 2820 1484
rect 2636 1376 2644 1384
rect 2556 1356 2564 1364
rect 2572 1356 2580 1364
rect 2620 1356 2628 1364
rect 2700 1396 2708 1404
rect 2748 1416 2756 1424
rect 2716 1376 2724 1384
rect 2748 1376 2756 1384
rect 2620 1336 2628 1344
rect 2668 1336 2676 1344
rect 2764 1336 2772 1344
rect 2492 1296 2500 1304
rect 2524 1296 2532 1304
rect 2380 1176 2388 1184
rect 2460 1176 2468 1184
rect 2460 1116 2468 1124
rect 2444 1056 2452 1064
rect 2428 1036 2436 1044
rect 2508 1196 2516 1204
rect 2604 1296 2612 1304
rect 2588 1256 2596 1264
rect 2572 1136 2580 1144
rect 2556 1096 2564 1104
rect 2524 1056 2532 1064
rect 2492 1016 2500 1024
rect 2380 956 2388 964
rect 2412 856 2420 864
rect 2428 856 2436 864
rect 2476 856 2484 864
rect 2492 796 2500 804
rect 2396 756 2404 764
rect 2444 756 2452 764
rect 2380 736 2388 744
rect 2332 676 2340 684
rect 2332 656 2340 664
rect 2284 516 2292 524
rect 2268 356 2276 364
rect 2252 296 2260 304
rect 2236 196 2244 204
rect 1852 136 1860 144
rect 1900 136 1908 144
rect 1964 136 1972 144
rect 2028 136 2036 144
rect 2140 136 2148 144
rect 1788 116 1796 124
rect 1868 116 1876 124
rect 1980 116 1988 124
rect 2108 116 2116 124
rect 2300 476 2308 484
rect 2412 716 2420 724
rect 2476 716 2484 724
rect 2492 716 2500 724
rect 2412 656 2420 664
rect 2364 516 2372 524
rect 2348 476 2356 484
rect 2348 416 2356 424
rect 2316 376 2324 384
rect 2444 576 2452 584
rect 2540 1016 2548 1024
rect 2540 936 2548 944
rect 2524 916 2532 924
rect 2524 796 2532 804
rect 2668 1316 2676 1324
rect 2748 1316 2756 1324
rect 2796 1316 2804 1324
rect 2812 1296 2820 1304
rect 2764 1256 2772 1264
rect 2860 1336 2868 1344
rect 3036 1796 3044 1804
rect 2988 1596 2996 1604
rect 2940 1556 2948 1564
rect 2956 1556 2964 1564
rect 2956 1536 2964 1544
rect 3148 1696 3156 1704
rect 3052 1536 3060 1544
rect 3004 1436 3012 1444
rect 2915 1406 2923 1414
rect 2925 1406 2933 1414
rect 2935 1406 2943 1414
rect 2945 1406 2953 1414
rect 2955 1406 2963 1414
rect 2965 1406 2973 1414
rect 2908 1336 2916 1344
rect 2860 1296 2868 1304
rect 2844 1236 2852 1244
rect 2620 1196 2628 1204
rect 2940 1296 2948 1304
rect 2908 1256 2916 1264
rect 2892 1116 2900 1124
rect 3020 1216 3028 1224
rect 3212 2036 3220 2044
rect 3276 1996 3284 2004
rect 3228 1976 3236 1984
rect 3180 1896 3188 1904
rect 3196 1876 3204 1884
rect 3180 1856 3188 1864
rect 3164 1616 3172 1624
rect 3164 1476 3172 1484
rect 3276 1956 3284 1964
rect 3244 1936 3252 1944
rect 3244 1896 3252 1904
rect 3260 1876 3268 1884
rect 3276 1836 3284 1844
rect 3260 1736 3268 1744
rect 3276 1736 3284 1744
rect 3196 1718 3204 1724
rect 3196 1716 3204 1718
rect 3244 1616 3252 1624
rect 3372 2136 3380 2144
rect 3436 2496 3444 2504
rect 3596 2796 3604 2804
rect 3644 2776 3652 2784
rect 3516 2756 3524 2764
rect 3548 2756 3556 2764
rect 3596 2756 3604 2764
rect 3676 2756 3684 2764
rect 3580 2736 3588 2744
rect 3500 2716 3508 2724
rect 3548 2716 3556 2724
rect 3676 2716 3684 2724
rect 3692 2716 3700 2724
rect 3596 2696 3604 2704
rect 3532 2656 3540 2664
rect 3564 2656 3572 2664
rect 3788 3056 3796 3064
rect 3820 3056 3828 3064
rect 3852 3056 3860 3064
rect 3788 3036 3796 3044
rect 3772 2996 3780 3004
rect 3836 3016 3844 3024
rect 3900 2996 3908 3004
rect 3788 2956 3796 2964
rect 3836 2956 3844 2964
rect 3740 2936 3748 2944
rect 3740 2896 3748 2904
rect 3964 3356 3972 3364
rect 4044 3476 4052 3484
rect 4012 3376 4020 3384
rect 4060 3356 4068 3364
rect 4044 3336 4052 3344
rect 3948 3316 3956 3324
rect 3996 3296 4004 3304
rect 4108 3336 4116 3344
rect 4092 3296 4100 3304
rect 4060 3276 4068 3284
rect 4028 3196 4036 3204
rect 3980 3116 3988 3124
rect 4252 3736 4260 3744
rect 4300 3776 4308 3784
rect 4492 4116 4500 4124
rect 4419 4006 4427 4014
rect 4429 4006 4437 4014
rect 4439 4006 4447 4014
rect 4449 4006 4457 4014
rect 4459 4006 4467 4014
rect 4469 4006 4477 4014
rect 4412 3902 4420 3904
rect 4412 3896 4420 3902
rect 4444 3896 4452 3904
rect 4476 3836 4484 3844
rect 4348 3796 4356 3804
rect 4412 3796 4420 3804
rect 4332 3736 4340 3744
rect 4348 3736 4356 3744
rect 4412 3736 4420 3744
rect 4220 3636 4228 3644
rect 4172 3536 4180 3544
rect 4172 3496 4180 3504
rect 4220 3496 4228 3504
rect 4284 3716 4292 3724
rect 4300 3696 4308 3704
rect 4300 3596 4308 3604
rect 4236 3356 4244 3364
rect 4284 3456 4292 3464
rect 4284 3376 4292 3384
rect 4252 3336 4260 3344
rect 4156 3316 4164 3324
rect 4380 3696 4388 3704
rect 4396 3676 4404 3684
rect 4380 3656 4388 3664
rect 4444 3656 4452 3664
rect 4364 3356 4372 3364
rect 4348 3336 4356 3344
rect 4332 3276 4340 3284
rect 4419 3606 4427 3614
rect 4429 3606 4437 3614
rect 4439 3606 4447 3614
rect 4449 3606 4457 3614
rect 4459 3606 4467 3614
rect 4469 3606 4477 3614
rect 4476 3576 4484 3584
rect 4412 3556 4420 3564
rect 4396 3496 4404 3504
rect 4412 3336 4420 3344
rect 4508 4016 4516 4024
rect 4572 4236 4580 4244
rect 4700 4496 4708 4504
rect 4796 4496 4804 4504
rect 4812 4496 4820 4504
rect 4844 4716 4852 4724
rect 5132 5036 5140 5044
rect 5116 4996 5124 5004
rect 5036 4856 5044 4864
rect 5084 4856 5092 4864
rect 4876 4716 4884 4724
rect 4956 4716 4964 4724
rect 5084 4716 5092 4724
rect 4956 4696 4964 4704
rect 4940 4676 4948 4684
rect 5132 4936 5140 4944
rect 5116 4916 5124 4924
rect 5116 4856 5124 4864
rect 5132 4756 5140 4764
rect 5212 5076 5220 5084
rect 5260 5056 5268 5064
rect 5308 5056 5316 5064
rect 5196 5036 5204 5044
rect 5180 4976 5188 4984
rect 5164 4956 5172 4964
rect 5212 4896 5220 4904
rect 5164 4756 5172 4764
rect 5148 4736 5156 4744
rect 5036 4676 5044 4684
rect 5004 4656 5012 4664
rect 4924 4636 4932 4644
rect 5068 4656 5076 4664
rect 5116 4656 5124 4664
rect 4860 4576 4868 4584
rect 4876 4576 4884 4584
rect 4844 4556 4852 4564
rect 4764 4476 4772 4484
rect 4812 4476 4820 4484
rect 4828 4476 4836 4484
rect 4764 4396 4772 4404
rect 4972 4616 4980 4624
rect 4940 4576 4948 4584
rect 4956 4556 4964 4564
rect 4892 4516 4900 4524
rect 4892 4496 4900 4504
rect 4812 4316 4820 4324
rect 4908 4476 4916 4484
rect 4796 4296 4804 4304
rect 4844 4296 4852 4304
rect 4652 4276 4660 4284
rect 4604 4236 4612 4244
rect 4636 4236 4644 4244
rect 4588 4196 4596 4204
rect 4892 4276 4900 4284
rect 4780 4236 4788 4244
rect 4732 4196 4740 4204
rect 4780 4196 4788 4204
rect 4716 4176 4724 4184
rect 4828 4176 4836 4184
rect 4876 4156 4884 4164
rect 4892 4156 4900 4164
rect 4748 4136 4756 4144
rect 4540 4116 4548 4124
rect 4604 4116 4612 4124
rect 4876 4116 4884 4124
rect 4780 4096 4788 4104
rect 4812 4096 4820 4104
rect 4860 4096 4868 4104
rect 4524 3996 4532 4004
rect 4652 3976 4660 3984
rect 4732 3976 4740 3984
rect 4508 3956 4516 3964
rect 4540 3836 4548 3844
rect 4604 3796 4612 3804
rect 4588 3776 4596 3784
rect 4524 3756 4532 3764
rect 4572 3736 4580 3744
rect 4556 3696 4564 3704
rect 4588 3716 4596 3724
rect 4668 3902 4676 3904
rect 4668 3896 4676 3902
rect 4700 3896 4708 3904
rect 4764 3836 4772 3844
rect 4700 3796 4708 3804
rect 4748 3796 4756 3804
rect 4796 3796 4804 3804
rect 4636 3736 4644 3744
rect 4668 3736 4676 3744
rect 4700 3736 4708 3744
rect 4780 3736 4788 3744
rect 4604 3676 4612 3684
rect 4572 3556 4580 3564
rect 4604 3456 4612 3464
rect 4492 3416 4500 3424
rect 4540 3436 4548 3444
rect 4540 3416 4548 3424
rect 4524 3396 4532 3404
rect 4508 3336 4516 3344
rect 4556 3396 4564 3404
rect 4572 3376 4580 3384
rect 4652 3576 4660 3584
rect 4668 3536 4676 3544
rect 4652 3496 4660 3504
rect 4732 3676 4740 3684
rect 4860 4076 4868 4084
rect 4860 3876 4868 3884
rect 4844 3856 4852 3864
rect 4956 4276 4964 4284
rect 4924 4176 4932 4184
rect 5020 4556 5028 4564
rect 5004 4456 5012 4464
rect 5052 4536 5060 4544
rect 5052 4516 5060 4524
rect 5036 4476 5044 4484
rect 5020 4396 5028 4404
rect 4988 4336 4996 4344
rect 5180 4716 5188 4724
rect 5212 4716 5220 4724
rect 5196 4596 5204 4604
rect 5308 4916 5316 4924
rect 5452 5236 5460 5244
rect 5404 5156 5412 5164
rect 5356 5136 5364 5144
rect 5372 5136 5380 5144
rect 5340 5056 5348 5064
rect 5436 5116 5444 5124
rect 5420 5096 5428 5104
rect 5404 5056 5412 5064
rect 5372 5036 5380 5044
rect 5436 5036 5444 5044
rect 5420 4976 5428 4984
rect 5356 4956 5364 4964
rect 5484 5176 5492 5184
rect 5500 5156 5508 5164
rect 5468 5076 5476 5084
rect 5660 5316 5668 5324
rect 5708 5316 5716 5324
rect 5628 5276 5636 5284
rect 5804 5356 5812 5364
rect 5900 5356 5908 5364
rect 5996 5356 6004 5364
rect 6188 5356 6196 5364
rect 6316 5356 6324 5364
rect 6412 5356 6420 5364
rect 6060 5336 6068 5344
rect 6124 5336 6132 5344
rect 6220 5336 6228 5344
rect 5772 5296 5780 5304
rect 5820 5296 5828 5304
rect 5852 5276 5860 5284
rect 5660 5216 5668 5224
rect 5724 5216 5732 5224
rect 5580 5176 5588 5184
rect 5548 5076 5556 5084
rect 5628 5076 5636 5084
rect 5516 4956 5524 4964
rect 5548 4956 5556 4964
rect 5420 4936 5428 4944
rect 5308 4816 5316 4824
rect 5468 4916 5476 4924
rect 5420 4756 5428 4764
rect 5372 4716 5380 4724
rect 5244 4656 5252 4664
rect 5324 4656 5332 4664
rect 5292 4636 5300 4644
rect 5260 4576 5268 4584
rect 5132 4556 5140 4564
rect 5228 4556 5236 4564
rect 5260 4556 5268 4564
rect 5084 4536 5092 4544
rect 5148 4536 5156 4544
rect 5244 4536 5252 4544
rect 5132 4516 5140 4524
rect 5212 4516 5220 4524
rect 5116 4496 5124 4504
rect 5068 4436 5076 4444
rect 5052 4396 5060 4404
rect 5068 4376 5076 4384
rect 5228 4476 5236 4484
rect 5148 4336 5156 4344
rect 5036 4296 5044 4304
rect 5084 4296 5092 4304
rect 5020 4256 5028 4264
rect 5004 4196 5012 4204
rect 4972 4156 4980 4164
rect 5020 4136 5028 4144
rect 4988 4116 4996 4124
rect 4956 4096 4964 4104
rect 5052 4096 5060 4104
rect 4908 4076 4916 4084
rect 4940 4076 4948 4084
rect 4908 4056 4916 4064
rect 4940 3936 4948 3944
rect 4908 3916 4916 3924
rect 4892 3816 4900 3824
rect 4892 3776 4900 3784
rect 4988 3916 4996 3924
rect 5020 3916 5028 3924
rect 4956 3896 4964 3904
rect 5212 4416 5220 4424
rect 5116 4276 5124 4284
rect 5132 4256 5140 4264
rect 5196 4256 5204 4264
rect 5148 4196 5156 4204
rect 5116 3936 5124 3944
rect 5084 3896 5092 3904
rect 5100 3896 5108 3904
rect 4956 3856 4964 3864
rect 4972 3856 4980 3864
rect 5036 3856 5044 3864
rect 4972 3816 4980 3824
rect 4972 3776 4980 3784
rect 5020 3776 5028 3784
rect 4876 3636 4884 3644
rect 4764 3616 4772 3624
rect 4812 3616 4820 3624
rect 4812 3536 4820 3544
rect 4764 3516 4772 3524
rect 4812 3516 4820 3524
rect 4828 3496 4836 3504
rect 4844 3496 4852 3504
rect 4732 3476 4740 3484
rect 4620 3416 4628 3424
rect 4684 3416 4692 3424
rect 4636 3336 4644 3344
rect 4524 3316 4532 3324
rect 4396 3296 4404 3304
rect 4476 3296 4484 3304
rect 4508 3296 4516 3304
rect 4419 3206 4427 3214
rect 4429 3206 4437 3214
rect 4439 3206 4447 3214
rect 4449 3206 4457 3214
rect 4459 3206 4467 3214
rect 4469 3206 4477 3214
rect 4204 3176 4212 3184
rect 4268 3176 4276 3184
rect 4284 3176 4292 3184
rect 4364 3176 4372 3184
rect 4380 3176 4388 3184
rect 4412 3176 4420 3184
rect 4156 3116 4164 3124
rect 4284 3116 4292 3124
rect 3996 3102 4004 3104
rect 3996 3096 4004 3102
rect 4124 3096 4132 3104
rect 4156 3096 4164 3104
rect 4220 3096 4228 3104
rect 4236 3096 4244 3104
rect 3980 3076 3988 3084
rect 4140 3076 4148 3084
rect 4172 3076 4180 3084
rect 4092 3056 4100 3064
rect 3980 3036 3988 3044
rect 4028 3016 4036 3024
rect 4076 3016 4084 3024
rect 3932 2936 3940 2944
rect 3996 2936 4004 2944
rect 3804 2916 3812 2924
rect 3964 2916 3972 2924
rect 3772 2796 3780 2804
rect 3756 2776 3764 2784
rect 3740 2756 3748 2764
rect 3724 2696 3732 2704
rect 3660 2656 3668 2664
rect 3644 2596 3652 2604
rect 3676 2636 3684 2644
rect 3564 2556 3572 2564
rect 3580 2556 3588 2564
rect 3644 2556 3652 2564
rect 3660 2556 3668 2564
rect 3628 2536 3636 2544
rect 3500 2518 3508 2524
rect 3500 2516 3508 2518
rect 3564 2516 3572 2524
rect 3628 2496 3636 2504
rect 3660 2536 3668 2544
rect 3676 2536 3684 2544
rect 3676 2496 3684 2504
rect 3484 2436 3492 2444
rect 3516 2436 3524 2444
rect 3596 2436 3604 2444
rect 3452 2416 3460 2424
rect 3468 2416 3476 2424
rect 3468 2356 3476 2364
rect 3500 2296 3508 2304
rect 3468 2256 3476 2264
rect 3404 2196 3412 2204
rect 3436 2196 3444 2204
rect 3452 2196 3460 2204
rect 3404 2176 3412 2184
rect 3452 2156 3460 2164
rect 3468 2156 3476 2164
rect 3708 2656 3716 2664
rect 3724 2656 3732 2664
rect 3900 2896 3908 2904
rect 3820 2876 3828 2884
rect 3884 2876 3892 2884
rect 3804 2736 3812 2744
rect 3868 2756 3876 2764
rect 3836 2736 3844 2744
rect 3836 2656 3844 2664
rect 3772 2576 3780 2584
rect 3788 2576 3796 2584
rect 3740 2556 3748 2564
rect 3756 2556 3764 2564
rect 3724 2516 3732 2524
rect 3692 2396 3700 2404
rect 3580 2356 3588 2364
rect 3596 2336 3604 2344
rect 3612 2316 3620 2324
rect 3644 2316 3652 2324
rect 3548 2296 3556 2304
rect 3596 2296 3604 2304
rect 3548 2276 3556 2284
rect 3532 2216 3540 2224
rect 3516 2156 3524 2164
rect 3468 2136 3476 2144
rect 3484 2136 3492 2144
rect 3500 2136 3508 2144
rect 3596 2236 3604 2244
rect 3564 2156 3572 2164
rect 3452 2056 3460 2064
rect 3372 2016 3380 2024
rect 3388 2016 3396 2024
rect 3340 1976 3348 1984
rect 3356 1976 3364 1984
rect 3340 1956 3348 1964
rect 3308 1896 3316 1904
rect 3324 1876 3332 1884
rect 3436 1996 3444 2004
rect 3356 1896 3364 1904
rect 3404 1876 3412 1884
rect 3356 1856 3364 1864
rect 3340 1796 3348 1804
rect 3388 1796 3396 1804
rect 3452 1896 3460 1904
rect 3468 1876 3476 1884
rect 3484 1876 3492 1884
rect 3468 1836 3476 1844
rect 3388 1776 3396 1784
rect 3452 1776 3460 1784
rect 3356 1736 3364 1744
rect 3372 1736 3380 1744
rect 3324 1676 3332 1684
rect 3324 1616 3332 1624
rect 3308 1516 3316 1524
rect 3196 1496 3204 1504
rect 3228 1496 3236 1504
rect 3244 1496 3252 1504
rect 3292 1496 3300 1504
rect 3372 1496 3380 1504
rect 3420 1496 3428 1504
rect 3212 1476 3220 1484
rect 3132 1436 3140 1444
rect 3180 1436 3188 1444
rect 3116 1416 3124 1424
rect 3148 1416 3156 1424
rect 3100 1356 3108 1364
rect 3100 1336 3108 1344
rect 3052 1156 3060 1164
rect 3100 1136 3108 1144
rect 2604 1056 2612 1064
rect 2572 736 2580 744
rect 2572 716 2580 724
rect 2556 696 2564 704
rect 2524 656 2532 664
rect 2556 656 2564 664
rect 2508 576 2516 584
rect 2428 556 2436 564
rect 2476 556 2484 564
rect 2620 1036 2628 1044
rect 2796 1102 2804 1104
rect 2796 1096 2804 1102
rect 2828 1096 2836 1104
rect 2908 1096 2916 1104
rect 3196 1396 3204 1404
rect 3148 1356 3156 1364
rect 3228 1356 3236 1364
rect 3212 1336 3220 1344
rect 3228 1336 3236 1344
rect 3148 1318 3156 1324
rect 3148 1316 3156 1318
rect 3292 1476 3300 1484
rect 3308 1476 3316 1484
rect 3356 1476 3364 1484
rect 3420 1476 3428 1484
rect 3436 1476 3444 1484
rect 3340 1436 3348 1444
rect 3388 1436 3396 1444
rect 3420 1436 3428 1444
rect 3372 1396 3380 1404
rect 3324 1336 3332 1344
rect 3276 1316 3284 1324
rect 3324 1316 3332 1324
rect 3260 1296 3268 1304
rect 3244 1256 3252 1264
rect 3244 1236 3252 1244
rect 3388 1236 3396 1244
rect 3228 1156 3236 1164
rect 3212 1096 3220 1104
rect 2876 1076 2884 1084
rect 3180 1076 3188 1084
rect 3212 1076 3220 1084
rect 2908 1056 2916 1064
rect 3276 1096 3284 1104
rect 3340 1096 3348 1104
rect 2636 996 2644 1004
rect 2636 956 2644 964
rect 2604 896 2612 904
rect 2620 856 2628 864
rect 2876 1016 2884 1024
rect 2988 1016 2996 1024
rect 2812 976 2820 984
rect 2844 936 2852 944
rect 2668 916 2676 924
rect 2915 1006 2923 1014
rect 2925 1006 2933 1014
rect 2935 1006 2943 1014
rect 2945 1006 2953 1014
rect 2955 1006 2963 1014
rect 2965 1006 2973 1014
rect 2892 996 2900 1004
rect 2652 836 2660 844
rect 2684 836 2692 844
rect 3244 1036 3252 1044
rect 3324 1036 3332 1044
rect 3164 976 3172 984
rect 3196 976 3204 984
rect 3116 936 3124 944
rect 3196 916 3204 924
rect 2748 816 2756 824
rect 2892 816 2900 824
rect 2684 776 2692 784
rect 2732 776 2740 784
rect 2620 716 2628 724
rect 2668 716 2676 724
rect 2428 536 2436 544
rect 2492 536 2500 544
rect 2396 496 2404 504
rect 2428 496 2436 504
rect 2380 336 2388 344
rect 2364 316 2372 324
rect 2364 296 2372 304
rect 2412 276 2420 284
rect 2412 236 2420 244
rect 2284 116 2292 124
rect 2348 196 2356 204
rect 2316 176 2324 184
rect 2508 516 2516 524
rect 2524 516 2532 524
rect 2476 496 2484 504
rect 2492 476 2500 484
rect 2460 396 2468 404
rect 2540 496 2548 504
rect 2636 656 2644 664
rect 2652 596 2660 604
rect 2588 556 2596 564
rect 2620 556 2628 564
rect 2652 536 2660 544
rect 2780 756 2788 764
rect 2828 736 2836 744
rect 2876 736 2884 744
rect 2892 736 2900 744
rect 2860 716 2868 724
rect 2732 636 2740 644
rect 2844 676 2852 684
rect 2748 616 2756 624
rect 2780 556 2788 564
rect 2796 536 2804 544
rect 2892 656 2900 664
rect 3036 876 3044 884
rect 3100 876 3108 884
rect 3020 776 3028 784
rect 2924 756 2932 764
rect 3020 736 3028 744
rect 2940 716 2948 724
rect 3068 716 3076 724
rect 3132 836 3140 844
rect 3036 676 3044 684
rect 3084 676 3092 684
rect 3004 656 3012 664
rect 3052 656 3060 664
rect 3196 816 3204 824
rect 3468 1736 3476 1744
rect 3500 1796 3508 1804
rect 3500 1776 3508 1784
rect 3548 2036 3556 2044
rect 3676 2296 3684 2304
rect 3724 2416 3732 2424
rect 3708 2356 3716 2364
rect 3628 2276 3636 2284
rect 3660 2256 3668 2264
rect 3628 2236 3636 2244
rect 3660 2216 3668 2224
rect 3692 2276 3700 2284
rect 3708 2276 3716 2284
rect 3612 2176 3620 2184
rect 3756 2496 3764 2504
rect 3756 2436 3764 2444
rect 3772 2436 3780 2444
rect 3772 2416 3780 2424
rect 3740 2336 3748 2344
rect 3932 2876 3940 2884
rect 3948 2856 3956 2864
rect 3900 2636 3908 2644
rect 3980 2776 3988 2784
rect 3964 2756 3972 2764
rect 4012 2916 4020 2924
rect 4316 3096 4324 3104
rect 4300 3056 4308 3064
rect 4204 3036 4212 3044
rect 4236 3036 4244 3044
rect 4172 2996 4180 3004
rect 4156 2976 4164 2984
rect 4076 2916 4084 2924
rect 4188 2936 4196 2944
rect 4124 2916 4132 2924
rect 4156 2916 4164 2924
rect 4092 2896 4100 2904
rect 4060 2876 4068 2884
rect 4044 2756 4052 2764
rect 4108 2876 4116 2884
rect 4172 2756 4180 2764
rect 4060 2736 4068 2744
rect 4092 2736 4100 2744
rect 4108 2736 4116 2744
rect 3996 2676 4004 2684
rect 3884 2596 3892 2604
rect 3916 2596 3924 2604
rect 3948 2596 3956 2604
rect 3868 2576 3876 2584
rect 3804 2556 3812 2564
rect 3836 2556 3844 2564
rect 3868 2556 3876 2564
rect 3820 2536 3828 2544
rect 3868 2516 3876 2524
rect 3916 2556 3924 2564
rect 3932 2556 3940 2564
rect 3868 2436 3876 2444
rect 3900 2416 3908 2424
rect 3820 2396 3828 2404
rect 3772 2316 3780 2324
rect 3756 2296 3764 2304
rect 3740 2236 3748 2244
rect 3580 2136 3588 2144
rect 3596 2136 3604 2144
rect 3580 2016 3588 2024
rect 3564 1956 3572 1964
rect 3548 1896 3556 1904
rect 3516 1736 3524 1744
rect 3548 1736 3556 1744
rect 3484 1716 3492 1724
rect 3468 1676 3476 1684
rect 3516 1676 3524 1684
rect 3644 2116 3652 2124
rect 3612 1896 3620 1904
rect 3772 2236 3780 2244
rect 3900 2336 3908 2344
rect 3868 2316 3876 2324
rect 3836 2276 3844 2284
rect 3852 2256 3860 2264
rect 3884 2276 3892 2284
rect 3868 2236 3876 2244
rect 3772 2176 3780 2184
rect 3836 2176 3844 2184
rect 3772 2116 3780 2124
rect 3788 2116 3796 2124
rect 3676 2036 3684 2044
rect 3724 2036 3732 2044
rect 3756 2036 3764 2044
rect 3628 1836 3636 1844
rect 3628 1816 3636 1824
rect 3612 1676 3620 1684
rect 3532 1516 3540 1524
rect 3548 1516 3556 1524
rect 3484 1496 3492 1504
rect 3548 1476 3556 1484
rect 3500 1436 3508 1444
rect 3468 1376 3476 1384
rect 3516 1356 3524 1364
rect 3580 1436 3588 1444
rect 3596 1436 3604 1444
rect 3596 1416 3604 1424
rect 3532 1336 3540 1344
rect 3564 1336 3572 1344
rect 3452 1316 3460 1324
rect 3468 1316 3476 1324
rect 3532 1316 3540 1324
rect 3692 1896 3700 1904
rect 3756 1996 3764 2004
rect 3676 1876 3684 1884
rect 3708 1876 3716 1884
rect 3740 1876 3748 1884
rect 3660 1836 3668 1844
rect 3676 1836 3684 1844
rect 3644 1776 3652 1784
rect 3676 1756 3684 1764
rect 3724 1756 3732 1764
rect 3836 2096 3844 2104
rect 3868 2096 3876 2104
rect 3804 2036 3812 2044
rect 3788 1996 3796 2004
rect 3852 1916 3860 1924
rect 3868 1896 3876 1904
rect 3804 1876 3812 1884
rect 3788 1836 3796 1844
rect 3868 1876 3876 1884
rect 3836 1856 3844 1864
rect 3820 1836 3828 1844
rect 3836 1796 3844 1804
rect 4012 2656 4020 2664
rect 3996 2636 4004 2644
rect 3980 2576 3988 2584
rect 3980 2556 3988 2564
rect 3964 2516 3972 2524
rect 4156 2716 4164 2724
rect 4188 2716 4196 2724
rect 4156 2696 4164 2704
rect 4172 2696 4180 2704
rect 4108 2656 4116 2664
rect 4140 2656 4148 2664
rect 4156 2656 4164 2664
rect 4204 2656 4212 2664
rect 4076 2596 4084 2604
rect 4092 2596 4100 2604
rect 4076 2576 4084 2584
rect 4028 2556 4036 2564
rect 4060 2556 4068 2564
rect 4028 2516 4036 2524
rect 4044 2516 4052 2524
rect 4124 2596 4132 2604
rect 4124 2576 4132 2584
rect 4092 2556 4100 2564
rect 4012 2476 4020 2484
rect 3964 2336 3972 2344
rect 3932 2316 3940 2324
rect 3996 2316 4004 2324
rect 4012 2316 4020 2324
rect 3980 2296 3988 2304
rect 3948 2276 3956 2284
rect 3964 2276 3972 2284
rect 3996 2256 4004 2264
rect 3948 2216 3956 2224
rect 3932 2196 3940 2204
rect 3932 2096 3940 2104
rect 3916 1896 3924 1904
rect 3900 1776 3908 1784
rect 3980 2176 3988 2184
rect 3996 2176 4004 2184
rect 3964 1996 3972 2004
rect 4092 2496 4100 2504
rect 4108 2496 4116 2504
rect 4044 2416 4052 2424
rect 4092 2416 4100 2424
rect 4188 2536 4196 2544
rect 4172 2516 4180 2524
rect 4300 2996 4308 3004
rect 4316 2936 4324 2944
rect 4348 3056 4356 3064
rect 4364 3036 4372 3044
rect 4492 3136 4500 3144
rect 4476 3096 4484 3104
rect 4572 3276 4580 3284
rect 4540 3176 4548 3184
rect 4412 3016 4420 3024
rect 4268 2916 4276 2924
rect 4284 2916 4292 2924
rect 4332 2916 4340 2924
rect 4364 2916 4372 2924
rect 4412 2976 4420 2984
rect 4316 2896 4324 2904
rect 4348 2876 4356 2884
rect 4252 2856 4260 2864
rect 4268 2856 4276 2864
rect 4236 2736 4244 2744
rect 4220 2596 4228 2604
rect 4332 2816 4340 2824
rect 4428 2916 4436 2924
rect 4412 2856 4420 2864
rect 4419 2806 4427 2814
rect 4429 2806 4437 2814
rect 4439 2806 4447 2814
rect 4449 2806 4457 2814
rect 4459 2806 4467 2814
rect 4469 2806 4477 2814
rect 4380 2796 4388 2804
rect 4540 3016 4548 3024
rect 4588 3096 4596 3104
rect 4620 3236 4628 3244
rect 4604 3016 4612 3024
rect 4604 2996 4612 3004
rect 4524 2956 4532 2964
rect 4540 2956 4548 2964
rect 4588 2956 4596 2964
rect 4508 2936 4516 2944
rect 4604 2876 4612 2884
rect 4588 2796 4596 2804
rect 4732 3436 4740 3444
rect 4828 3396 4836 3404
rect 4764 3376 4772 3384
rect 4860 3376 4868 3384
rect 4700 3336 4708 3344
rect 4796 3336 4804 3344
rect 4844 3316 4852 3324
rect 4844 3296 4852 3304
rect 4732 3196 4740 3204
rect 4780 3196 4788 3204
rect 4716 3096 4724 3104
rect 4940 3736 4948 3744
rect 4924 3716 4932 3724
rect 5084 3816 5092 3824
rect 5068 3796 5076 3804
rect 5084 3796 5092 3804
rect 5116 3796 5124 3804
rect 5052 3756 5060 3764
rect 5036 3736 5044 3744
rect 5004 3716 5012 3724
rect 4988 3656 4996 3664
rect 4924 3476 4932 3484
rect 4924 3436 4932 3444
rect 4908 3396 4916 3404
rect 4876 3236 4884 3244
rect 4636 2956 4644 2964
rect 4668 2816 4676 2824
rect 4412 2776 4420 2784
rect 4364 2716 4372 2724
rect 4252 2656 4260 2664
rect 4252 2596 4260 2604
rect 4220 2496 4228 2504
rect 4204 2416 4212 2424
rect 4220 2416 4228 2424
rect 4076 2336 4084 2344
rect 4044 2296 4052 2304
rect 4188 2376 4196 2384
rect 4204 2376 4212 2384
rect 4124 2356 4132 2364
rect 4108 2276 4116 2284
rect 4172 2276 4180 2284
rect 4156 2256 4164 2264
rect 4060 2236 4068 2244
rect 4076 2236 4084 2244
rect 4028 2216 4036 2224
rect 4204 2256 4212 2264
rect 4188 2236 4196 2244
rect 4108 2196 4116 2204
rect 4156 2216 4164 2224
rect 4092 2156 4100 2164
rect 4124 2156 4132 2164
rect 4252 2476 4260 2484
rect 4252 2436 4260 2444
rect 4236 2396 4244 2404
rect 4252 2396 4260 2404
rect 4252 2356 4260 2364
rect 4300 2656 4308 2664
rect 4284 2616 4292 2624
rect 4284 2576 4292 2584
rect 4332 2516 4340 2524
rect 4748 3016 4756 3024
rect 4812 2976 4820 2984
rect 4748 2856 4756 2864
rect 4652 2756 4660 2764
rect 4684 2756 4692 2764
rect 4492 2736 4500 2744
rect 4556 2736 4564 2744
rect 4284 2436 4292 2444
rect 4268 2296 4276 2304
rect 4236 2216 4244 2224
rect 4188 2156 4196 2164
rect 4252 2156 4260 2164
rect 4028 2116 4036 2124
rect 4140 2116 4148 2124
rect 4236 2116 4244 2124
rect 4252 2116 4260 2124
rect 4012 2096 4020 2104
rect 4044 2096 4052 2104
rect 4204 2096 4212 2104
rect 4012 2076 4020 2084
rect 4028 2076 4036 2084
rect 4060 2076 4068 2084
rect 4028 2036 4036 2044
rect 3964 1916 3972 1924
rect 4060 1996 4068 2004
rect 4124 1996 4132 2004
rect 4076 1916 4084 1924
rect 4108 1916 4116 1924
rect 3980 1876 3988 1884
rect 4044 1876 4052 1884
rect 3932 1856 3940 1864
rect 3980 1856 3988 1864
rect 3996 1856 4004 1864
rect 4044 1856 4052 1864
rect 4076 1856 4084 1864
rect 4012 1816 4020 1824
rect 4028 1776 4036 1784
rect 3916 1756 3924 1764
rect 4012 1756 4020 1764
rect 4060 1756 4068 1764
rect 4172 1956 4180 1964
rect 4188 1956 4196 1964
rect 4220 2016 4228 2024
rect 4236 2016 4244 2024
rect 4252 1996 4260 2004
rect 4220 1916 4228 1924
rect 4140 1876 4148 1884
rect 4204 1876 4212 1884
rect 4188 1856 4196 1864
rect 3900 1736 3908 1744
rect 3964 1736 3972 1744
rect 3804 1716 3812 1724
rect 3644 1676 3652 1684
rect 3676 1676 3684 1684
rect 3692 1676 3700 1684
rect 3644 1616 3652 1624
rect 3644 1476 3652 1484
rect 3628 1416 3636 1424
rect 3628 1356 3636 1364
rect 3436 1296 3444 1304
rect 3564 1296 3572 1304
rect 3564 1256 3572 1264
rect 3500 1196 3508 1204
rect 3548 1196 3556 1204
rect 3484 1116 3492 1124
rect 3404 976 3412 984
rect 3420 976 3428 984
rect 3356 936 3364 944
rect 3388 916 3396 924
rect 3468 1096 3476 1104
rect 3532 1096 3540 1104
rect 3468 1076 3476 1084
rect 3548 1076 3556 1084
rect 3452 1056 3460 1064
rect 3500 1056 3508 1064
rect 3516 1036 3524 1044
rect 3500 996 3508 1004
rect 3484 976 3492 984
rect 3468 956 3476 964
rect 3452 936 3460 944
rect 3484 936 3492 944
rect 3516 936 3524 944
rect 3532 876 3540 884
rect 3612 1316 3620 1324
rect 3724 1636 3732 1644
rect 3708 1616 3716 1624
rect 3676 1476 3684 1484
rect 3708 1476 3716 1484
rect 3660 1436 3668 1444
rect 3676 1416 3684 1424
rect 3708 1416 3716 1424
rect 3788 1656 3796 1664
rect 3772 1616 3780 1624
rect 3740 1496 3748 1504
rect 3772 1496 3780 1504
rect 3804 1556 3812 1564
rect 3932 1716 3940 1724
rect 3884 1616 3892 1624
rect 3900 1616 3908 1624
rect 3836 1596 3844 1604
rect 3900 1576 3908 1584
rect 3868 1516 3876 1524
rect 3756 1436 3764 1444
rect 3788 1476 3796 1484
rect 3724 1316 3732 1324
rect 3660 1296 3668 1304
rect 3580 1016 3588 1024
rect 3596 1016 3604 1024
rect 3644 996 3652 1004
rect 3740 1256 3748 1264
rect 3692 1116 3700 1124
rect 3772 1396 3780 1404
rect 3788 1276 3796 1284
rect 3692 1102 3700 1104
rect 3692 1096 3700 1102
rect 3756 1096 3764 1104
rect 3612 936 3620 944
rect 3820 1476 3828 1484
rect 3868 1456 3876 1464
rect 3948 1596 3956 1604
rect 3996 1636 4004 1644
rect 4076 1736 4084 1744
rect 3932 1576 3940 1584
rect 3948 1576 3956 1584
rect 3916 1496 3924 1504
rect 3852 1436 3860 1444
rect 3916 1456 3924 1464
rect 3900 1416 3908 1424
rect 3996 1536 4004 1544
rect 3980 1436 3988 1444
rect 3964 1356 3972 1364
rect 3948 1336 3956 1344
rect 3852 1296 3860 1304
rect 3868 1296 3876 1304
rect 3852 1276 3860 1284
rect 3836 1256 3844 1264
rect 3836 1216 3844 1224
rect 3724 996 3732 1004
rect 3772 1016 3780 1024
rect 3692 936 3700 944
rect 3756 936 3764 944
rect 3804 976 3812 984
rect 3852 1176 3860 1184
rect 3916 1296 3924 1304
rect 3884 1116 3892 1124
rect 3868 1036 3876 1044
rect 3868 1016 3876 1024
rect 3788 936 3796 944
rect 3820 936 3828 944
rect 3676 916 3684 924
rect 3564 836 3572 844
rect 3516 776 3524 784
rect 3500 756 3508 764
rect 3148 676 3156 684
rect 2908 636 2916 644
rect 3052 636 3060 644
rect 2915 606 2923 614
rect 2925 606 2933 614
rect 2935 606 2943 614
rect 2945 606 2953 614
rect 2955 606 2963 614
rect 2965 606 2973 614
rect 2924 576 2932 584
rect 2844 556 2852 564
rect 2908 556 2916 564
rect 2716 516 2724 524
rect 2748 516 2756 524
rect 2812 516 2820 524
rect 2636 496 2644 504
rect 2572 396 2580 404
rect 2508 376 2516 384
rect 2636 416 2644 424
rect 2668 376 2676 384
rect 2620 356 2628 364
rect 2604 336 2612 344
rect 2636 336 2644 344
rect 2508 296 2516 304
rect 2444 256 2452 264
rect 2428 216 2436 224
rect 2476 256 2484 264
rect 2540 276 2548 284
rect 2540 256 2548 264
rect 2684 276 2692 284
rect 2524 236 2532 244
rect 2588 236 2596 244
rect 2492 176 2500 184
rect 2396 136 2404 144
rect 2476 136 2484 144
rect 2588 196 2596 204
rect 2812 356 2820 364
rect 2716 336 2724 344
rect 2732 296 2740 304
rect 2764 296 2772 304
rect 2700 256 2708 264
rect 2796 256 2804 264
rect 2764 236 2772 244
rect 2844 296 2852 304
rect 2844 256 2852 264
rect 2876 516 2884 524
rect 2908 476 2916 484
rect 2908 316 2916 324
rect 3036 556 3044 564
rect 3020 536 3028 544
rect 2956 296 2964 304
rect 2988 276 2996 284
rect 2876 216 2884 224
rect 2915 206 2923 214
rect 2925 206 2933 214
rect 2935 206 2943 214
rect 2945 206 2953 214
rect 2955 206 2963 214
rect 2965 206 2973 214
rect 2860 196 2868 204
rect 2716 176 2724 184
rect 2764 176 2772 184
rect 2812 176 2820 184
rect 2604 156 2612 164
rect 2668 156 2676 164
rect 2732 156 2740 164
rect 2620 136 2628 144
rect 2636 136 2644 144
rect 2780 136 2788 144
rect 3132 536 3140 544
rect 3052 396 3060 404
rect 3164 496 3172 504
rect 3132 376 3140 384
rect 3164 376 3172 384
rect 3116 356 3124 364
rect 3100 336 3108 344
rect 3068 316 3076 324
rect 3132 316 3140 324
rect 3116 296 3124 304
rect 3068 256 3076 264
rect 3036 176 3044 184
rect 3116 176 3124 184
rect 3052 156 3060 164
rect 2908 136 2916 144
rect 3004 136 3012 144
rect 3148 296 3156 304
rect 3148 276 3156 284
rect 3404 696 3412 704
rect 3484 696 3492 704
rect 3388 676 3396 684
rect 3260 536 3268 544
rect 3420 536 3428 544
rect 3484 596 3492 604
rect 3596 816 3604 824
rect 3644 816 3652 824
rect 3580 536 3588 544
rect 3292 518 3300 524
rect 3292 516 3300 518
rect 3468 516 3476 524
rect 3708 856 3716 864
rect 3756 896 3764 904
rect 3724 836 3732 844
rect 3756 816 3764 824
rect 3724 696 3732 704
rect 3612 576 3620 584
rect 3676 496 3684 504
rect 3356 396 3364 404
rect 3500 376 3508 384
rect 3548 376 3556 384
rect 3372 356 3380 364
rect 3340 336 3348 344
rect 3292 296 3300 304
rect 3228 276 3236 284
rect 3276 276 3284 284
rect 3228 256 3236 264
rect 3148 236 3156 244
rect 3196 136 3204 144
rect 3244 196 3252 204
rect 3404 276 3412 284
rect 3372 176 3380 184
rect 3340 156 3348 164
rect 2348 116 2356 124
rect 2652 116 2660 124
rect 2684 116 2692 124
rect 2764 116 2772 124
rect 2796 116 2804 124
rect 3660 316 3668 324
rect 3532 302 3540 304
rect 3532 296 3540 302
rect 3660 156 3668 164
rect 3740 518 3748 524
rect 3740 516 3748 518
rect 3836 896 3844 904
rect 4140 1756 4148 1764
rect 4188 1756 4196 1764
rect 4316 2296 4324 2304
rect 4300 2236 4308 2244
rect 4316 2236 4324 2244
rect 4284 2176 4292 2184
rect 4460 2496 4468 2504
rect 4412 2456 4420 2464
rect 4419 2406 4427 2414
rect 4429 2406 4437 2414
rect 4439 2406 4447 2414
rect 4449 2406 4457 2414
rect 4459 2406 4467 2414
rect 4469 2406 4477 2414
rect 4396 2396 4404 2404
rect 4604 2716 4612 2724
rect 4540 2656 4548 2664
rect 4556 2656 4564 2664
rect 4508 2576 4516 2584
rect 4540 2556 4548 2564
rect 4524 2536 4532 2544
rect 4508 2516 4516 2524
rect 4508 2496 4516 2504
rect 4492 2356 4500 2364
rect 4492 2336 4500 2344
rect 4428 2316 4436 2324
rect 4396 2296 4404 2304
rect 4332 2216 4340 2224
rect 4364 2156 4372 2164
rect 4348 2116 4356 2124
rect 4316 2076 4324 2084
rect 4348 2096 4356 2104
rect 4364 2096 4372 2104
rect 4284 1956 4292 1964
rect 4332 1956 4340 1964
rect 4268 1876 4276 1884
rect 4252 1856 4260 1864
rect 4300 1856 4308 1864
rect 4236 1776 4244 1784
rect 4124 1736 4132 1744
rect 4172 1736 4180 1744
rect 4124 1716 4132 1724
rect 4156 1656 4164 1664
rect 4108 1556 4116 1564
rect 4108 1536 4116 1544
rect 4012 1496 4020 1504
rect 4092 1476 4100 1484
rect 4044 1456 4052 1464
rect 4076 1456 4084 1464
rect 4028 1436 4036 1444
rect 4092 1436 4100 1444
rect 4044 1376 4052 1384
rect 3996 1356 4004 1364
rect 4012 1356 4020 1364
rect 4012 1336 4020 1344
rect 3996 1316 4004 1324
rect 3980 1296 3988 1304
rect 3964 1276 3972 1284
rect 3980 1236 3988 1244
rect 3932 1216 3940 1224
rect 4012 1176 4020 1184
rect 4124 1496 4132 1504
rect 4076 1356 4084 1364
rect 4044 1336 4052 1344
rect 4044 1296 4052 1304
rect 4076 1296 4084 1304
rect 4060 1276 4068 1284
rect 4076 1276 4084 1284
rect 3948 1136 3956 1144
rect 3980 1136 3988 1144
rect 3996 1136 4004 1144
rect 3932 1096 3940 1104
rect 3964 1096 3972 1104
rect 3980 1096 3988 1104
rect 3932 1076 3940 1084
rect 3884 956 3892 964
rect 3916 996 3924 1004
rect 4028 1116 4036 1124
rect 4044 1096 4052 1104
rect 4012 1076 4020 1084
rect 3932 976 3940 984
rect 3916 956 3924 964
rect 3932 936 3940 944
rect 3964 936 3972 944
rect 3868 896 3876 904
rect 3868 856 3876 864
rect 3868 816 3876 824
rect 3804 716 3812 724
rect 3932 716 3940 724
rect 3948 716 3956 724
rect 3804 696 3812 704
rect 4060 1076 4068 1084
rect 4060 1056 4068 1064
rect 4028 996 4036 1004
rect 4012 896 4020 904
rect 3980 816 3988 824
rect 4012 776 4020 784
rect 3980 736 3988 744
rect 3916 696 3924 704
rect 3964 696 3972 704
rect 3948 676 3956 684
rect 4044 976 4052 984
rect 4044 956 4052 964
rect 4108 1276 4116 1284
rect 4108 1256 4116 1264
rect 4092 1176 4100 1184
rect 4204 1656 4212 1664
rect 4204 1476 4212 1484
rect 4188 1456 4196 1464
rect 4188 1416 4196 1424
rect 4140 1316 4148 1324
rect 4156 1316 4164 1324
rect 4092 1136 4100 1144
rect 4108 1116 4116 1124
rect 4108 996 4116 1004
rect 4236 1756 4244 1764
rect 4396 2096 4404 2104
rect 4524 2476 4532 2484
rect 4524 2456 4532 2464
rect 4572 2596 4580 2604
rect 4588 2556 4596 2564
rect 4572 2516 4580 2524
rect 4540 2396 4548 2404
rect 4636 2676 4644 2684
rect 4636 2616 4644 2624
rect 4620 2576 4628 2584
rect 4604 2496 4612 2504
rect 4684 2576 4692 2584
rect 4716 2616 4724 2624
rect 4844 2776 4852 2784
rect 4844 2696 4852 2704
rect 4780 2676 4788 2684
rect 4716 2576 4724 2584
rect 4732 2576 4740 2584
rect 4700 2556 4708 2564
rect 4652 2536 4660 2544
rect 4700 2536 4708 2544
rect 4732 2536 4740 2544
rect 4684 2516 4692 2524
rect 4636 2476 4644 2484
rect 4668 2416 4676 2424
rect 4540 2356 4548 2364
rect 4556 2356 4564 2364
rect 4620 2356 4628 2364
rect 4636 2356 4644 2364
rect 4652 2316 4660 2324
rect 4556 2276 4564 2284
rect 4636 2276 4644 2284
rect 4732 2516 4740 2524
rect 4716 2396 4724 2404
rect 4700 2376 4708 2384
rect 4716 2316 4724 2324
rect 4700 2296 4708 2304
rect 4828 2616 4836 2624
rect 4764 2576 4772 2584
rect 4780 2576 4788 2584
rect 4812 2556 4820 2564
rect 4780 2536 4788 2544
rect 4764 2516 4772 2524
rect 4748 2316 4756 2324
rect 4748 2296 4756 2304
rect 4732 2256 4740 2264
rect 4572 2236 4580 2244
rect 4684 2236 4692 2244
rect 4508 2156 4516 2164
rect 4540 2136 4548 2144
rect 4492 2116 4500 2124
rect 4476 2096 4484 2104
rect 4412 2076 4420 2084
rect 4380 2016 4388 2024
rect 4419 2006 4427 2014
rect 4429 2006 4437 2014
rect 4439 2006 4447 2014
rect 4449 2006 4457 2014
rect 4459 2006 4467 2014
rect 4469 2006 4477 2014
rect 4380 1976 4388 1984
rect 4396 1976 4404 1984
rect 4444 1976 4452 1984
rect 4460 1976 4468 1984
rect 4428 1916 4436 1924
rect 4364 1896 4372 1904
rect 4364 1816 4372 1824
rect 4364 1776 4372 1784
rect 4236 1476 4244 1484
rect 4236 1456 4244 1464
rect 4220 1276 4228 1284
rect 4172 1236 4180 1244
rect 4156 1196 4164 1204
rect 4156 1156 4164 1164
rect 4140 1056 4148 1064
rect 4092 976 4100 984
rect 4124 976 4132 984
rect 4092 896 4100 904
rect 4124 896 4132 904
rect 4316 1736 4324 1744
rect 4380 1656 4388 1664
rect 4508 2036 4516 2044
rect 4748 2216 4756 2224
rect 4620 2196 4628 2204
rect 4588 2140 4596 2144
rect 4588 2136 4596 2140
rect 4604 2136 4612 2144
rect 4780 2436 4788 2444
rect 4812 2316 4820 2324
rect 4796 2256 4804 2264
rect 4828 2196 4836 2204
rect 4668 2176 4676 2184
rect 4876 2976 4884 2984
rect 4972 3396 4980 3404
rect 4956 3356 4964 3364
rect 5020 3456 5028 3464
rect 5180 4176 5188 4184
rect 5308 4516 5316 4524
rect 5292 4496 5300 4504
rect 5308 4456 5316 4464
rect 5260 4336 5268 4344
rect 5228 4156 5236 4164
rect 5228 4136 5236 4144
rect 5324 4416 5332 4424
rect 5356 4596 5364 4604
rect 5484 4756 5492 4764
rect 5452 4696 5460 4704
rect 5644 4956 5652 4964
rect 5596 4896 5604 4904
rect 5564 4856 5572 4864
rect 5580 4856 5588 4864
rect 5596 4816 5604 4824
rect 5580 4776 5588 4784
rect 5596 4776 5604 4784
rect 5564 4756 5572 4764
rect 5500 4616 5508 4624
rect 5548 4616 5556 4624
rect 5388 4596 5396 4604
rect 5484 4596 5492 4604
rect 5436 4576 5444 4584
rect 5532 4596 5540 4604
rect 5804 5136 5812 5144
rect 5724 5116 5732 5124
rect 5676 5056 5684 5064
rect 5724 5056 5732 5064
rect 5740 5036 5748 5044
rect 5708 5016 5716 5024
rect 5692 4996 5700 5004
rect 5692 4956 5700 4964
rect 5724 4936 5732 4944
rect 5756 4936 5764 4944
rect 5836 5116 5844 5124
rect 5900 5256 5908 5264
rect 5884 5136 5892 5144
rect 5868 5116 5876 5124
rect 5884 5096 5892 5104
rect 5820 5076 5828 5084
rect 5804 5036 5812 5044
rect 5852 5036 5860 5044
rect 5788 5016 5796 5024
rect 6124 5196 6132 5204
rect 6364 5336 6372 5344
rect 6460 5336 6468 5344
rect 6796 5336 6804 5344
rect 6220 5316 6228 5324
rect 6268 5316 6276 5324
rect 6364 5296 6372 5304
rect 6284 5216 6292 5224
rect 5996 5156 6004 5164
rect 6156 5156 6164 5164
rect 5916 5096 5924 5104
rect 6012 5136 6020 5144
rect 6156 5136 6164 5144
rect 6220 5116 6228 5124
rect 6172 5096 6180 5104
rect 6188 5096 6196 5104
rect 6028 5056 6036 5064
rect 6108 5056 6116 5064
rect 6332 5176 6340 5184
rect 6332 5156 6340 5164
rect 6300 5116 6308 5124
rect 6268 5096 6276 5104
rect 6268 5076 6276 5084
rect 6220 5056 6228 5064
rect 6252 5056 6260 5064
rect 5932 5036 5940 5044
rect 6172 5036 6180 5044
rect 6268 5036 6276 5044
rect 5900 5016 5908 5024
rect 5923 5006 5931 5014
rect 5933 5006 5941 5014
rect 5943 5006 5951 5014
rect 5953 5006 5961 5014
rect 5963 5006 5971 5014
rect 5973 5006 5981 5014
rect 5852 4996 5860 5004
rect 6076 4996 6084 5004
rect 5804 4936 5812 4944
rect 5724 4916 5732 4924
rect 5740 4916 5748 4924
rect 5772 4916 5780 4924
rect 5692 4856 5700 4864
rect 5660 4756 5668 4764
rect 5708 4696 5716 4704
rect 5788 4896 5796 4904
rect 5756 4856 5764 4864
rect 5756 4836 5764 4844
rect 5788 4836 5796 4844
rect 5740 4736 5748 4744
rect 5628 4676 5636 4684
rect 5884 4976 5892 4984
rect 6012 4956 6020 4964
rect 6188 4976 6196 4984
rect 6140 4956 6148 4964
rect 6204 4956 6212 4964
rect 6172 4936 6180 4944
rect 5852 4916 5860 4924
rect 5964 4916 5972 4924
rect 6028 4916 6036 4924
rect 5788 4756 5796 4764
rect 5804 4756 5812 4764
rect 5772 4736 5780 4744
rect 5580 4556 5588 4564
rect 5724 4656 5732 4664
rect 5740 4656 5748 4664
rect 5628 4636 5636 4644
rect 5660 4636 5668 4644
rect 5388 4516 5396 4524
rect 5468 4516 5476 4524
rect 5596 4516 5604 4524
rect 5612 4516 5620 4524
rect 5356 4496 5364 4504
rect 5500 4456 5508 4464
rect 5404 4416 5412 4424
rect 5436 4356 5444 4364
rect 5340 4336 5348 4344
rect 5564 4336 5572 4344
rect 5484 4296 5492 4304
rect 5308 4276 5316 4284
rect 5340 4276 5348 4284
rect 5292 4236 5300 4244
rect 5276 4156 5284 4164
rect 5292 4156 5300 4164
rect 5244 4096 5252 4104
rect 5260 4036 5268 4044
rect 5244 3976 5252 3984
rect 5212 3916 5220 3924
rect 5196 3896 5204 3904
rect 5180 3816 5188 3824
rect 5164 3796 5172 3804
rect 5228 3856 5236 3864
rect 5260 3936 5268 3944
rect 5324 4256 5332 4264
rect 5340 4256 5348 4264
rect 5420 4256 5428 4264
rect 5372 4236 5380 4244
rect 5532 4276 5540 4284
rect 5564 4256 5572 4264
rect 5500 4236 5508 4244
rect 5548 4236 5556 4244
rect 5612 4336 5620 4344
rect 5612 4296 5620 4304
rect 5596 4256 5604 4264
rect 5468 4216 5476 4224
rect 5356 4196 5364 4204
rect 5388 4196 5396 4204
rect 5308 4096 5316 4104
rect 5388 4096 5396 4104
rect 5292 4076 5300 4084
rect 5404 4076 5412 4084
rect 5292 3936 5300 3944
rect 5484 3936 5492 3944
rect 5324 3916 5332 3924
rect 5212 3836 5220 3844
rect 5244 3836 5252 3844
rect 5148 3756 5156 3764
rect 5196 3756 5204 3764
rect 5100 3716 5108 3724
rect 5276 3856 5284 3864
rect 5228 3816 5236 3824
rect 5260 3816 5268 3824
rect 5276 3816 5284 3824
rect 5164 3736 5172 3744
rect 5116 3696 5124 3704
rect 5084 3656 5092 3664
rect 5116 3496 5124 3504
rect 5100 3476 5108 3484
rect 5132 3476 5140 3484
rect 5004 3376 5012 3384
rect 5036 3376 5044 3384
rect 5084 3376 5092 3384
rect 5276 3756 5284 3764
rect 5180 3716 5188 3724
rect 5244 3716 5252 3724
rect 5276 3696 5284 3704
rect 5532 4196 5540 4204
rect 5516 4056 5524 4064
rect 5564 4176 5572 4184
rect 5612 4236 5620 4244
rect 5612 4196 5620 4204
rect 5612 4156 5620 4164
rect 5532 3976 5540 3984
rect 5612 4116 5620 4124
rect 5612 4056 5620 4064
rect 5596 3916 5604 3924
rect 5500 3896 5508 3904
rect 5420 3876 5428 3884
rect 5452 3856 5460 3864
rect 5484 3836 5492 3844
rect 5340 3816 5348 3824
rect 5420 3796 5428 3804
rect 5324 3736 5332 3744
rect 5468 3736 5476 3744
rect 5356 3676 5364 3684
rect 5292 3656 5300 3664
rect 5532 3876 5540 3884
rect 5516 3816 5524 3824
rect 5564 3816 5572 3824
rect 5596 3776 5604 3784
rect 5452 3716 5460 3724
rect 5500 3716 5508 3724
rect 5532 3716 5540 3724
rect 5404 3696 5412 3704
rect 5420 3696 5428 3704
rect 5420 3556 5428 3564
rect 5228 3496 5236 3504
rect 5260 3502 5268 3504
rect 5260 3496 5268 3502
rect 5292 3496 5300 3504
rect 5436 3496 5444 3504
rect 5180 3396 5188 3404
rect 5068 3356 5076 3364
rect 5148 3356 5156 3364
rect 5004 3316 5012 3324
rect 5148 3316 5156 3324
rect 5292 3416 5300 3424
rect 5388 3476 5396 3484
rect 5404 3456 5412 3464
rect 5420 3396 5428 3404
rect 5340 3376 5348 3384
rect 5372 3376 5380 3384
rect 5212 3336 5220 3344
rect 5404 3336 5412 3344
rect 5244 3318 5252 3324
rect 5244 3316 5252 3318
rect 5116 3276 5124 3284
rect 5164 3276 5172 3284
rect 5244 3276 5252 3284
rect 4988 3256 4996 3264
rect 5036 3256 5044 3264
rect 5132 3256 5140 3264
rect 5068 3116 5076 3124
rect 5148 3116 5156 3124
rect 5228 3116 5236 3124
rect 4940 3096 4948 3104
rect 5068 3096 5076 3104
rect 5180 3096 5188 3104
rect 5196 3096 5204 3104
rect 5052 3036 5060 3044
rect 4892 2936 4900 2944
rect 4892 2916 4900 2924
rect 4876 2696 4884 2704
rect 4876 2596 4884 2604
rect 5100 2996 5108 3004
rect 5020 2956 5028 2964
rect 5052 2936 5060 2944
rect 5164 3056 5172 3064
rect 5164 3036 5172 3044
rect 5196 2976 5204 2984
rect 5212 2976 5220 2984
rect 5516 3696 5524 3704
rect 5724 4616 5732 4624
rect 5692 4596 5700 4604
rect 5660 4576 5668 4584
rect 5676 4556 5684 4564
rect 5836 4896 5844 4904
rect 5820 4716 5828 4724
rect 5788 4656 5796 4664
rect 5820 4576 5828 4584
rect 5756 4556 5764 4564
rect 5868 4876 5876 4884
rect 6092 4856 6100 4864
rect 6156 4876 6164 4884
rect 6044 4816 6052 4824
rect 6108 4816 6116 4824
rect 5916 4796 5924 4804
rect 6140 4796 6148 4804
rect 5868 4756 5876 4764
rect 5900 4756 5908 4764
rect 6108 4756 6116 4764
rect 5964 4716 5972 4724
rect 6060 4716 6068 4724
rect 5948 4696 5956 4704
rect 5996 4696 6004 4704
rect 6012 4676 6020 4684
rect 5996 4616 6004 4624
rect 5923 4606 5931 4614
rect 5933 4606 5941 4614
rect 5943 4606 5951 4614
rect 5953 4606 5961 4614
rect 5963 4606 5971 4614
rect 5973 4606 5981 4614
rect 5900 4596 5908 4604
rect 5692 4536 5700 4544
rect 5708 4536 5716 4544
rect 5644 4516 5652 4524
rect 5804 4496 5812 4504
rect 5660 4456 5668 4464
rect 5644 4316 5652 4324
rect 5644 4256 5652 4264
rect 5820 4416 5828 4424
rect 5836 4416 5844 4424
rect 5804 4376 5812 4384
rect 5708 4336 5716 4344
rect 5676 4316 5684 4324
rect 5820 4316 5828 4324
rect 5756 4296 5764 4304
rect 5772 4296 5780 4304
rect 5804 4296 5812 4304
rect 5708 4276 5716 4284
rect 5740 4276 5748 4284
rect 5724 4256 5732 4264
rect 5724 4236 5732 4244
rect 5660 4156 5668 4164
rect 5756 4196 5764 4204
rect 5724 4136 5732 4144
rect 5692 4096 5700 4104
rect 5772 4156 5780 4164
rect 5772 4136 5780 4144
rect 5868 4536 5876 4544
rect 6044 4596 6052 4604
rect 5980 4536 5988 4544
rect 5900 4496 5908 4504
rect 5884 4296 5892 4304
rect 6220 4936 6228 4944
rect 6284 4996 6292 5004
rect 6348 4996 6356 5004
rect 6524 5296 6532 5304
rect 6572 5296 6580 5304
rect 6476 5276 6484 5284
rect 6540 5276 6548 5284
rect 6572 5276 6580 5284
rect 6428 5256 6436 5264
rect 6460 5116 6468 5124
rect 6524 5076 6532 5084
rect 6412 5056 6420 5064
rect 6492 5036 6500 5044
rect 6460 5016 6468 5024
rect 6396 4976 6404 4984
rect 6428 4976 6436 4984
rect 6332 4936 6340 4944
rect 6364 4936 6372 4944
rect 6460 4956 6468 4964
rect 6444 4936 6452 4944
rect 6524 4976 6532 4984
rect 6572 5236 6580 5244
rect 6556 5096 6564 5104
rect 6716 5276 6724 5284
rect 6588 5216 6596 5224
rect 6636 5116 6644 5124
rect 6988 5376 6996 5384
rect 7196 5356 7204 5364
rect 7068 5336 7076 5344
rect 6716 5096 6724 5104
rect 6764 5096 6772 5104
rect 6828 5096 6836 5104
rect 6572 5076 6580 5084
rect 6556 4996 6564 5004
rect 7020 5316 7028 5324
rect 7164 5316 7172 5324
rect 7308 5316 7316 5324
rect 7004 5236 7012 5244
rect 6988 5136 6996 5144
rect 6636 5076 6644 5084
rect 6908 5076 6916 5084
rect 6956 5076 6964 5084
rect 6604 5036 6612 5044
rect 6796 4996 6804 5004
rect 6588 4956 6596 4964
rect 6940 4976 6948 4984
rect 6652 4956 6660 4964
rect 6908 4956 6916 4964
rect 6988 4956 6996 4964
rect 6668 4936 6676 4944
rect 6684 4936 6692 4944
rect 6780 4936 6788 4944
rect 6268 4876 6276 4884
rect 6300 4916 6308 4924
rect 6380 4916 6388 4924
rect 6476 4916 6484 4924
rect 6300 4856 6308 4864
rect 6412 4856 6420 4864
rect 6204 4836 6212 4844
rect 6284 4836 6292 4844
rect 6076 4696 6084 4704
rect 6124 4696 6132 4704
rect 6156 4696 6164 4704
rect 6092 4656 6100 4664
rect 6044 4496 6052 4504
rect 6060 4496 6068 4504
rect 6028 4456 6036 4464
rect 5884 4276 5892 4284
rect 5916 4276 5924 4284
rect 5868 4256 5876 4264
rect 5852 4236 5860 4244
rect 5852 4216 5860 4224
rect 5836 4196 5844 4204
rect 5884 4156 5892 4164
rect 5923 4206 5931 4214
rect 5933 4206 5941 4214
rect 5943 4206 5951 4214
rect 5953 4206 5961 4214
rect 5963 4206 5971 4214
rect 5973 4206 5981 4214
rect 5884 4136 5892 4144
rect 5884 4116 5892 4124
rect 5660 4076 5668 4084
rect 5708 4076 5716 4084
rect 5788 4076 5796 4084
rect 5788 4036 5796 4044
rect 5932 4156 5940 4164
rect 5948 4116 5956 4124
rect 5724 3976 5732 3984
rect 5788 3976 5796 3984
rect 5916 3976 5924 3984
rect 5660 3936 5668 3944
rect 5772 3936 5780 3944
rect 5692 3856 5700 3864
rect 5756 3856 5764 3864
rect 5644 3776 5652 3784
rect 5644 3736 5652 3744
rect 5628 3676 5636 3684
rect 5644 3656 5652 3664
rect 5580 3636 5588 3644
rect 5580 3576 5588 3584
rect 5580 3536 5588 3544
rect 5516 3496 5524 3504
rect 5484 3476 5492 3484
rect 5532 3476 5540 3484
rect 5452 3456 5460 3464
rect 5452 3416 5460 3424
rect 5452 3316 5460 3324
rect 5436 3196 5444 3204
rect 5324 3136 5332 3144
rect 5388 3136 5396 3144
rect 5340 3096 5348 3104
rect 5452 3096 5460 3104
rect 5260 2996 5268 3004
rect 5292 2976 5300 2984
rect 5308 2976 5316 2984
rect 5228 2936 5236 2944
rect 5244 2916 5252 2924
rect 5020 2856 5028 2864
rect 5228 2896 5236 2904
rect 5228 2856 5236 2864
rect 5340 2936 5348 2944
rect 5324 2916 5332 2924
rect 5340 2896 5348 2904
rect 5308 2836 5316 2844
rect 5324 2776 5332 2784
rect 5100 2736 5108 2744
rect 5068 2716 5076 2724
rect 5004 2696 5012 2704
rect 4956 2676 4964 2684
rect 4924 2636 4932 2644
rect 4956 2636 4964 2644
rect 4908 2516 4916 2524
rect 4940 2616 4948 2624
rect 5020 2616 5028 2624
rect 4940 2576 4948 2584
rect 5004 2556 5012 2564
rect 4860 2496 4868 2504
rect 4860 2456 4868 2464
rect 4716 2136 4724 2144
rect 4636 2116 4644 2124
rect 4604 2096 4612 2104
rect 4572 1976 4580 1984
rect 4540 1956 4548 1964
rect 4604 1956 4612 1964
rect 4524 1896 4532 1904
rect 4492 1876 4500 1884
rect 4588 1916 4596 1924
rect 4524 1856 4532 1864
rect 4556 1856 4564 1864
rect 4492 1776 4500 1784
rect 4460 1756 4468 1764
rect 4524 1756 4532 1764
rect 4572 1756 4580 1764
rect 4540 1736 4548 1744
rect 4460 1716 4468 1724
rect 4476 1716 4484 1724
rect 4508 1696 4516 1704
rect 4524 1696 4532 1704
rect 4348 1636 4356 1644
rect 4380 1636 4388 1644
rect 4396 1636 4404 1644
rect 4444 1636 4452 1644
rect 4460 1636 4468 1644
rect 4268 1576 4276 1584
rect 4364 1576 4372 1584
rect 4332 1536 4340 1544
rect 4300 1516 4308 1524
rect 4252 1416 4260 1424
rect 4252 1356 4260 1364
rect 4268 1296 4276 1304
rect 4252 1136 4260 1144
rect 4316 1236 4324 1244
rect 4284 1176 4292 1184
rect 4204 1096 4212 1104
rect 4268 1096 4276 1104
rect 4172 1076 4180 1084
rect 4188 1076 4196 1084
rect 4188 1036 4196 1044
rect 4156 776 4164 784
rect 4044 716 4052 724
rect 4076 716 4084 724
rect 3836 636 3844 644
rect 3820 616 3828 624
rect 3788 596 3796 604
rect 3820 556 3828 564
rect 3900 656 3908 664
rect 3996 656 4004 664
rect 4028 656 4036 664
rect 3900 596 3908 604
rect 4044 596 4052 604
rect 3980 576 3988 584
rect 3868 556 3876 564
rect 3916 556 3924 564
rect 3980 556 3988 564
rect 4044 556 4052 564
rect 4076 556 4084 564
rect 3804 516 3812 524
rect 3868 516 3876 524
rect 3948 536 3956 544
rect 3964 536 3972 544
rect 4012 516 4020 524
rect 3932 496 3940 504
rect 4012 496 4020 504
rect 3772 396 3780 404
rect 3852 396 3860 404
rect 3772 376 3780 384
rect 3948 356 3956 364
rect 3868 316 3876 324
rect 3884 316 3892 324
rect 3932 296 3940 304
rect 3756 256 3764 264
rect 3788 256 3796 264
rect 3804 256 3812 264
rect 3836 236 3844 244
rect 3868 256 3876 264
rect 3852 196 3860 204
rect 3820 176 3828 184
rect 3852 176 3860 184
rect 3724 156 3732 164
rect 3708 136 3716 144
rect 3836 136 3844 144
rect 3932 236 3940 244
rect 3932 196 3940 204
rect 4076 518 4084 524
rect 4076 516 4084 518
rect 4124 736 4132 744
rect 4156 736 4164 744
rect 4284 1076 4292 1084
rect 4236 996 4244 1004
rect 4252 976 4260 984
rect 4284 956 4292 964
rect 4419 1606 4427 1614
rect 4429 1606 4437 1614
rect 4439 1606 4447 1614
rect 4449 1606 4457 1614
rect 4459 1606 4467 1614
rect 4469 1606 4477 1614
rect 4492 1596 4500 1604
rect 4556 1656 4564 1664
rect 4540 1636 4548 1644
rect 4348 1496 4356 1504
rect 4348 1296 4356 1304
rect 4364 1296 4372 1304
rect 4492 1556 4500 1564
rect 4508 1556 4516 1564
rect 4396 1536 4404 1544
rect 4412 1496 4420 1504
rect 4508 1456 4516 1464
rect 4524 1456 4532 1464
rect 4444 1376 4452 1384
rect 4524 1376 4532 1384
rect 4508 1356 4516 1364
rect 4348 1216 4356 1224
rect 4332 1136 4340 1144
rect 4348 1136 4356 1144
rect 4348 1116 4356 1124
rect 4332 1096 4340 1104
rect 4316 936 4324 944
rect 4348 916 4356 924
rect 4316 896 4324 904
rect 4380 1096 4388 1104
rect 4220 816 4228 824
rect 4252 816 4260 824
rect 4236 776 4244 784
rect 4364 856 4372 864
rect 4188 756 4196 764
rect 4236 756 4244 764
rect 4268 756 4276 764
rect 4220 716 4228 724
rect 4284 716 4292 724
rect 4172 696 4180 704
rect 4252 696 4260 704
rect 4108 676 4116 684
rect 4172 676 4180 684
rect 4220 676 4228 684
rect 4188 656 4196 664
rect 4156 636 4164 644
rect 4108 616 4116 624
rect 4204 616 4212 624
rect 4428 1236 4436 1244
rect 4492 1216 4500 1224
rect 4419 1206 4427 1214
rect 4429 1206 4437 1214
rect 4439 1206 4447 1214
rect 4449 1206 4457 1214
rect 4459 1206 4467 1214
rect 4469 1206 4477 1214
rect 4428 1176 4436 1184
rect 4476 1176 4484 1184
rect 4508 1196 4516 1204
rect 4492 1136 4500 1144
rect 4604 1876 4612 1884
rect 4620 1856 4628 1864
rect 4620 1736 4628 1744
rect 4604 1716 4612 1724
rect 4620 1716 4628 1724
rect 4588 1516 4596 1524
rect 4572 1476 4580 1484
rect 4556 1416 4564 1424
rect 4588 1416 4596 1424
rect 4540 1256 4548 1264
rect 4540 1236 4548 1244
rect 4524 1176 4532 1184
rect 4444 1096 4452 1104
rect 4508 1096 4516 1104
rect 4412 976 4420 984
rect 4620 1676 4628 1684
rect 4716 2116 4724 2124
rect 4700 2036 4708 2044
rect 4700 1876 4708 1884
rect 4764 2096 4772 2104
rect 4796 2096 4804 2104
rect 4780 2056 4788 2064
rect 4908 2416 4916 2424
rect 4956 2216 4964 2224
rect 4940 2176 4948 2184
rect 4876 2136 4884 2144
rect 4876 2036 4884 2044
rect 4908 2036 4916 2044
rect 4828 1956 4836 1964
rect 4732 1936 4740 1944
rect 4764 1916 4772 1924
rect 4716 1856 4724 1864
rect 4684 1756 4692 1764
rect 4668 1736 4676 1744
rect 4716 1736 4724 1744
rect 4716 1676 4724 1684
rect 4684 1636 4692 1644
rect 4652 1536 4660 1544
rect 4636 1496 4644 1504
rect 4620 1476 4628 1484
rect 4604 1276 4612 1284
rect 4620 1256 4628 1264
rect 4700 1556 4708 1564
rect 4748 1856 4756 1864
rect 4780 1736 4788 1744
rect 4780 1716 4788 1724
rect 4764 1656 4772 1664
rect 4844 1896 4852 1904
rect 4892 1876 4900 1884
rect 4844 1796 4852 1804
rect 4972 2016 4980 2024
rect 5148 2716 5156 2724
rect 5228 2716 5236 2724
rect 5148 2696 5156 2704
rect 5164 2696 5172 2704
rect 5196 2696 5204 2704
rect 5212 2656 5220 2664
rect 5196 2616 5204 2624
rect 5132 2456 5140 2464
rect 5100 2356 5108 2364
rect 5052 2336 5060 2344
rect 5052 2296 5060 2304
rect 5068 2296 5076 2304
rect 5116 2296 5124 2304
rect 5148 2356 5156 2364
rect 5052 2276 5060 2284
rect 5084 2276 5092 2284
rect 5068 2236 5076 2244
rect 5148 2236 5156 2244
rect 5116 2216 5124 2224
rect 5004 2136 5012 2144
rect 5004 2116 5012 2124
rect 5052 2116 5060 2124
rect 5228 2516 5236 2524
rect 5196 2396 5204 2404
rect 5196 2336 5204 2344
rect 5212 2296 5220 2304
rect 5228 2296 5236 2304
rect 5180 2276 5188 2284
rect 5180 2196 5188 2204
rect 5276 2576 5284 2584
rect 5372 3076 5380 3084
rect 5436 3036 5444 3044
rect 5356 2876 5364 2884
rect 5452 2996 5460 3004
rect 5564 3416 5572 3424
rect 5612 3476 5620 3484
rect 5644 3476 5652 3484
rect 5628 3436 5636 3444
rect 5596 3356 5604 3364
rect 5612 3316 5620 3324
rect 5564 3296 5572 3304
rect 5532 3276 5540 3284
rect 5564 3276 5572 3284
rect 5692 3836 5700 3844
rect 5756 3816 5764 3824
rect 5756 3776 5764 3784
rect 5740 3736 5748 3744
rect 5676 3716 5684 3724
rect 5676 3596 5684 3604
rect 5724 3716 5732 3724
rect 5692 3556 5700 3564
rect 5708 3556 5716 3564
rect 5884 3916 5892 3924
rect 5836 3896 5844 3904
rect 5820 3876 5828 3884
rect 5804 3856 5812 3864
rect 5836 3696 5844 3704
rect 5836 3676 5844 3684
rect 5788 3536 5796 3544
rect 5708 3496 5716 3504
rect 5756 3496 5764 3504
rect 5788 3496 5796 3504
rect 5820 3496 5828 3504
rect 5692 3436 5700 3444
rect 5804 3476 5812 3484
rect 5724 3376 5732 3384
rect 5660 3276 5668 3284
rect 5676 3276 5684 3284
rect 5596 3256 5604 3264
rect 5644 3256 5652 3264
rect 5676 3256 5684 3264
rect 5644 3196 5652 3204
rect 5788 3356 5796 3364
rect 5756 3336 5764 3344
rect 5724 3296 5732 3304
rect 5708 3256 5716 3264
rect 5692 3216 5700 3224
rect 5612 3156 5620 3164
rect 5516 3116 5524 3124
rect 5564 3096 5572 3104
rect 5500 3076 5508 3084
rect 5484 3036 5492 3044
rect 5580 3036 5588 3044
rect 5404 2936 5412 2944
rect 5500 2936 5508 2944
rect 5436 2916 5444 2924
rect 5404 2896 5412 2904
rect 5388 2776 5396 2784
rect 5436 2756 5444 2764
rect 5340 2696 5348 2704
rect 5484 2736 5492 2744
rect 5500 2696 5508 2704
rect 5404 2676 5412 2684
rect 5468 2676 5476 2684
rect 5372 2656 5380 2664
rect 5436 2656 5444 2664
rect 5484 2656 5492 2664
rect 5372 2616 5380 2624
rect 5452 2556 5460 2564
rect 5308 2516 5316 2524
rect 5276 2376 5284 2384
rect 5404 2496 5412 2504
rect 5340 2476 5348 2484
rect 5388 2476 5396 2484
rect 5404 2456 5412 2464
rect 5420 2456 5428 2464
rect 5324 2416 5332 2424
rect 5308 2316 5316 2324
rect 5292 2276 5300 2284
rect 5164 2116 5172 2124
rect 5180 2116 5188 2124
rect 5260 2116 5268 2124
rect 5100 2056 5108 2064
rect 5148 2056 5156 2064
rect 5068 2036 5076 2044
rect 4988 1996 4996 2004
rect 5052 1996 5060 2004
rect 5004 1916 5012 1924
rect 5068 1976 5076 1984
rect 5132 1936 5140 1944
rect 5148 1916 5156 1924
rect 5244 2076 5252 2084
rect 5260 2076 5268 2084
rect 5292 2076 5300 2084
rect 5212 1916 5220 1924
rect 5020 1876 5028 1884
rect 5132 1876 5140 1884
rect 4924 1756 4932 1764
rect 4828 1736 4836 1744
rect 4876 1576 4884 1584
rect 4732 1516 4740 1524
rect 4668 1176 4676 1184
rect 4588 1136 4596 1144
rect 4652 1136 4660 1144
rect 4684 1156 4692 1164
rect 4604 1116 4612 1124
rect 4588 1096 4596 1104
rect 4652 1096 4660 1104
rect 4764 1536 4772 1544
rect 4828 1536 4836 1544
rect 4860 1516 4868 1524
rect 4780 1496 4788 1504
rect 4844 1496 4852 1504
rect 4796 1416 4804 1424
rect 4812 1376 4820 1384
rect 4748 1356 4756 1364
rect 4812 1356 4820 1364
rect 4828 1256 4836 1264
rect 4796 1176 4804 1184
rect 4732 1136 4740 1144
rect 4828 1136 4836 1144
rect 4748 1096 4756 1104
rect 4700 1076 4708 1084
rect 4572 1056 4580 1064
rect 4620 1056 4628 1064
rect 4524 1036 4532 1044
rect 4668 976 4676 984
rect 4684 976 4692 984
rect 4652 956 4660 964
rect 4540 936 4548 944
rect 4508 916 4516 924
rect 4572 896 4580 904
rect 4540 876 4548 884
rect 4604 856 4612 864
rect 4524 836 4532 844
rect 4540 836 4548 844
rect 4492 816 4500 824
rect 4419 806 4427 814
rect 4429 806 4437 814
rect 4439 806 4447 814
rect 4449 806 4457 814
rect 4459 806 4467 814
rect 4469 806 4477 814
rect 4396 776 4404 784
rect 4412 756 4420 764
rect 4140 516 4148 524
rect 4284 516 4292 524
rect 4220 476 4228 484
rect 4124 396 4132 404
rect 4092 376 4100 384
rect 4092 356 4100 364
rect 4156 356 4164 364
rect 4220 356 4228 364
rect 3996 316 4004 324
rect 4044 296 4052 304
rect 4028 276 4036 284
rect 3964 256 3972 264
rect 4044 256 4052 264
rect 4060 256 4068 264
rect 4028 236 4036 244
rect 4012 196 4020 204
rect 3916 156 3924 164
rect 3964 156 3972 164
rect 3996 156 4004 164
rect 4044 156 4052 164
rect 1772 96 1780 104
rect 1932 96 1940 104
rect 2300 96 2308 104
rect 3628 116 3636 124
rect 4092 256 4100 264
rect 4092 216 4100 224
rect 4076 176 4084 184
rect 4124 316 4132 324
rect 4172 316 4180 324
rect 4316 496 4324 504
rect 4748 936 4756 944
rect 4748 916 4756 924
rect 4908 1736 4916 1744
rect 4940 1736 4948 1744
rect 4940 1676 4948 1684
rect 4924 1636 4932 1644
rect 4924 1536 4932 1544
rect 4892 1476 4900 1484
rect 4860 1356 4868 1364
rect 4860 1136 4868 1144
rect 4860 1116 4868 1124
rect 5132 1856 5140 1864
rect 5116 1836 5124 1844
rect 5068 1756 5076 1764
rect 5036 1736 5044 1744
rect 4988 1716 4996 1724
rect 4972 1596 4980 1604
rect 5196 1536 5204 1544
rect 5004 1516 5012 1524
rect 5116 1516 5124 1524
rect 4956 1476 4964 1484
rect 4988 1416 4996 1424
rect 4908 1356 4916 1364
rect 4924 1356 4932 1364
rect 4908 1296 4916 1304
rect 4988 1296 4996 1304
rect 4924 1196 4932 1204
rect 4844 1096 4852 1104
rect 4892 1096 4900 1104
rect 4844 1076 4852 1084
rect 4780 1056 4788 1064
rect 4828 1056 4836 1064
rect 4780 1036 4788 1044
rect 4716 896 4724 904
rect 4700 796 4708 804
rect 4508 776 4516 784
rect 4524 776 4532 784
rect 4716 736 4724 744
rect 4764 896 4772 904
rect 4636 716 4644 724
rect 4748 716 4756 724
rect 4732 696 4740 704
rect 4540 676 4548 684
rect 4700 676 4708 684
rect 4492 596 4500 604
rect 4524 576 4532 584
rect 4652 596 4660 604
rect 4380 476 4388 484
rect 4419 406 4427 414
rect 4429 406 4437 414
rect 4439 406 4447 414
rect 4449 406 4457 414
rect 4459 406 4467 414
rect 4469 406 4477 414
rect 4332 396 4340 404
rect 4476 356 4484 364
rect 4204 276 4212 284
rect 4156 256 4164 264
rect 4172 216 4180 224
rect 4172 196 4180 204
rect 4252 156 4260 164
rect 4268 136 4276 144
rect 4380 276 4388 284
rect 4332 256 4340 264
rect 4380 256 4388 264
rect 4380 196 4388 204
rect 4492 196 4500 204
rect 4364 176 4372 184
rect 4396 156 4404 164
rect 4412 136 4420 144
rect 4540 276 4548 284
rect 4716 576 4724 584
rect 4716 516 4724 524
rect 4684 456 4692 464
rect 4748 556 4756 564
rect 4668 376 4676 384
rect 4700 316 4708 324
rect 4700 296 4708 304
rect 4748 296 4756 304
rect 4796 916 4804 924
rect 4796 856 4804 864
rect 4812 856 4820 864
rect 4812 776 4820 784
rect 4796 736 4804 744
rect 4812 736 4820 744
rect 4780 716 4788 724
rect 4812 676 4820 684
rect 4780 656 4788 664
rect 4812 616 4820 624
rect 4796 596 4804 604
rect 4812 556 4820 564
rect 4812 516 4820 524
rect 4780 496 4788 504
rect 4860 956 4868 964
rect 4860 936 4868 944
rect 4860 876 4868 884
rect 4844 796 4852 804
rect 4844 716 4852 724
rect 4892 976 4900 984
rect 4924 956 4932 964
rect 4892 936 4900 944
rect 4908 916 4916 924
rect 4892 776 4900 784
rect 4876 676 4884 684
rect 4844 656 4852 664
rect 4860 616 4868 624
rect 4876 556 4884 564
rect 4860 536 4868 544
rect 4860 516 4868 524
rect 4844 496 4852 504
rect 4828 356 4836 364
rect 4796 336 4804 344
rect 4812 336 4820 344
rect 4588 236 4596 244
rect 4716 236 4724 244
rect 4556 156 4564 164
rect 4508 116 4516 124
rect 3756 96 3764 104
rect 3996 96 4004 104
rect 4060 96 4068 104
rect 396 76 404 84
rect 460 76 468 84
rect 1276 76 1284 84
rect 1468 76 1476 84
rect 2284 76 2292 84
rect 2316 76 2324 84
rect 1411 6 1419 14
rect 1421 6 1429 14
rect 1431 6 1439 14
rect 1441 6 1449 14
rect 1451 6 1459 14
rect 1461 6 1469 14
rect 3500 16 3508 24
rect 3564 16 3572 24
rect 3660 16 3668 24
rect 4060 16 4068 24
rect 4419 6 4427 14
rect 4429 6 4437 14
rect 4439 6 4447 14
rect 4449 6 4457 14
rect 4459 6 4467 14
rect 4469 6 4477 14
rect 4572 136 4580 144
rect 4636 136 4644 144
rect 4700 136 4708 144
rect 4604 116 4612 124
rect 4652 116 4660 124
rect 4684 116 4692 124
rect 4748 156 4756 164
rect 4764 156 4772 164
rect 4588 96 4596 104
rect 4796 256 4804 264
rect 4796 216 4804 224
rect 4988 896 4996 904
rect 5100 1496 5108 1504
rect 5084 1436 5092 1444
rect 5164 1436 5172 1444
rect 5132 1416 5140 1424
rect 5100 1356 5108 1364
rect 5084 1316 5092 1324
rect 5164 1316 5172 1324
rect 5020 1136 5028 1144
rect 5228 1836 5236 1844
rect 5244 1796 5252 1804
rect 5276 1916 5284 1924
rect 5276 1736 5284 1744
rect 5404 2396 5412 2404
rect 5372 2376 5380 2384
rect 5372 2316 5380 2324
rect 5324 2296 5332 2304
rect 5340 2296 5348 2304
rect 5388 2296 5396 2304
rect 5324 2136 5332 2144
rect 5356 2276 5364 2284
rect 5420 2376 5428 2384
rect 5372 2216 5380 2224
rect 5356 2116 5364 2124
rect 5324 2036 5332 2044
rect 5308 1896 5316 1904
rect 5340 2016 5348 2024
rect 5404 2136 5412 2144
rect 5628 3036 5636 3044
rect 5644 2956 5652 2964
rect 5612 2836 5620 2844
rect 5596 2816 5604 2824
rect 5580 2736 5588 2744
rect 5548 2696 5556 2704
rect 5548 2676 5556 2684
rect 5516 2596 5524 2604
rect 5516 2556 5524 2564
rect 5532 2556 5540 2564
rect 5548 2536 5556 2544
rect 5564 2496 5572 2504
rect 5500 2456 5508 2464
rect 5596 2456 5604 2464
rect 5484 2416 5492 2424
rect 5580 2416 5588 2424
rect 5468 2316 5476 2324
rect 5500 2316 5508 2324
rect 5500 2276 5508 2284
rect 5500 2256 5508 2264
rect 5532 2256 5540 2264
rect 5436 2236 5444 2244
rect 5468 2236 5476 2244
rect 5484 2116 5492 2124
rect 5340 1976 5348 1984
rect 5372 1976 5380 1984
rect 5388 1976 5396 1984
rect 5308 1856 5316 1864
rect 5388 1816 5396 1824
rect 5372 1736 5380 1744
rect 5292 1716 5300 1724
rect 5228 1556 5236 1564
rect 5212 1516 5220 1524
rect 5292 1656 5300 1664
rect 5324 1716 5332 1724
rect 5340 1716 5348 1724
rect 5420 1996 5428 2004
rect 5420 1756 5428 1764
rect 5404 1676 5412 1684
rect 5420 1616 5428 1624
rect 5276 1576 5284 1584
rect 5404 1556 5412 1564
rect 5420 1556 5428 1564
rect 5388 1516 5396 1524
rect 5404 1516 5412 1524
rect 5308 1496 5316 1504
rect 5324 1496 5332 1504
rect 5372 1496 5380 1504
rect 5276 1476 5284 1484
rect 5292 1476 5300 1484
rect 5260 1416 5268 1424
rect 5244 1396 5252 1404
rect 5212 1376 5220 1384
rect 5308 1436 5316 1444
rect 5276 1356 5284 1364
rect 5196 1276 5204 1284
rect 5100 1256 5108 1264
rect 5116 1256 5124 1264
rect 5068 1176 5076 1184
rect 5052 1076 5060 1084
rect 5180 1176 5188 1184
rect 5132 1136 5140 1144
rect 5244 1136 5252 1144
rect 5132 1116 5140 1124
rect 5132 1076 5140 1084
rect 5100 1056 5108 1064
rect 5116 1016 5124 1024
rect 5100 956 5108 964
rect 5020 916 5028 924
rect 5036 896 5044 904
rect 5004 796 5012 804
rect 5212 1036 5220 1044
rect 5228 976 5236 984
rect 5212 956 5220 964
rect 5180 936 5188 944
rect 5164 916 5172 924
rect 5148 896 5156 904
rect 5132 876 5140 884
rect 5180 876 5188 884
rect 5516 2096 5524 2104
rect 5484 2036 5492 2044
rect 5564 2296 5572 2304
rect 5580 2256 5588 2264
rect 5580 2156 5588 2164
rect 5580 2116 5588 2124
rect 5564 2096 5572 2104
rect 5644 2816 5652 2824
rect 5724 3076 5732 3084
rect 5724 2796 5732 2804
rect 5708 2716 5716 2724
rect 5708 2696 5716 2704
rect 5644 2676 5652 2684
rect 5980 3896 5988 3904
rect 5948 3876 5956 3884
rect 5884 3836 5892 3844
rect 5923 3806 5931 3814
rect 5933 3806 5941 3814
rect 5943 3806 5951 3814
rect 5953 3806 5961 3814
rect 5963 3806 5971 3814
rect 5973 3806 5981 3814
rect 5900 3796 5908 3804
rect 5948 3776 5956 3784
rect 5964 3776 5972 3784
rect 6044 4256 6052 4264
rect 6012 4216 6020 4224
rect 6028 4176 6036 4184
rect 6092 4456 6100 4464
rect 6268 4776 6276 4784
rect 6380 4756 6388 4764
rect 6332 4716 6340 4724
rect 6348 4716 6356 4724
rect 6252 4696 6260 4704
rect 6204 4676 6212 4684
rect 6220 4676 6228 4684
rect 6172 4656 6180 4664
rect 6300 4656 6308 4664
rect 6140 4616 6148 4624
rect 6236 4616 6244 4624
rect 6268 4576 6276 4584
rect 6140 4536 6148 4544
rect 6204 4516 6212 4524
rect 6236 4516 6244 4524
rect 6172 4456 6180 4464
rect 6252 4436 6260 4444
rect 6108 4416 6116 4424
rect 6156 4416 6164 4424
rect 6092 4376 6100 4384
rect 6076 4316 6084 4324
rect 6236 4356 6244 4364
rect 6300 4516 6308 4524
rect 6284 4496 6292 4504
rect 6284 4456 6292 4464
rect 6172 4316 6180 4324
rect 6236 4316 6244 4324
rect 6268 4316 6276 4324
rect 6220 4256 6228 4264
rect 6076 4156 6084 4164
rect 6044 4116 6052 4124
rect 6092 4116 6100 4124
rect 6028 4076 6036 4084
rect 6044 4076 6052 4084
rect 6092 4056 6100 4064
rect 6044 4016 6052 4024
rect 6060 4016 6068 4024
rect 6044 3996 6052 4004
rect 6028 3956 6036 3964
rect 6044 3956 6052 3964
rect 6220 4236 6228 4244
rect 6220 4216 6228 4224
rect 6204 4196 6212 4204
rect 6156 4156 6164 4164
rect 6220 4156 6228 4164
rect 6124 4116 6132 4124
rect 6124 3996 6132 4004
rect 6108 3936 6116 3944
rect 6060 3916 6068 3924
rect 6012 3816 6020 3824
rect 6108 3856 6116 3864
rect 6076 3816 6084 3824
rect 6060 3796 6068 3804
rect 5868 3736 5876 3744
rect 6028 3776 6036 3784
rect 6108 3776 6116 3784
rect 6060 3736 6068 3744
rect 6092 3736 6100 3744
rect 6044 3716 6052 3724
rect 6012 3696 6020 3704
rect 6028 3696 6036 3704
rect 6028 3656 6036 3664
rect 6044 3656 6052 3664
rect 5980 3596 5988 3604
rect 6012 3596 6020 3604
rect 6076 3676 6084 3684
rect 6076 3656 6084 3664
rect 6060 3556 6068 3564
rect 6060 3516 6068 3524
rect 5996 3496 6004 3504
rect 6028 3496 6036 3504
rect 6044 3496 6052 3504
rect 5964 3456 5972 3464
rect 5900 3416 5908 3424
rect 5923 3406 5931 3414
rect 5933 3406 5941 3414
rect 5943 3406 5951 3414
rect 5953 3406 5961 3414
rect 5963 3406 5971 3414
rect 5973 3406 5981 3414
rect 5836 3256 5844 3264
rect 5820 3156 5828 3164
rect 5820 3116 5828 3124
rect 5756 3096 5764 3104
rect 5772 3096 5780 3104
rect 5804 3096 5812 3104
rect 6172 4116 6180 4124
rect 6156 3956 6164 3964
rect 6140 3916 6148 3924
rect 6188 4056 6196 4064
rect 6220 3996 6228 4004
rect 6188 3956 6196 3964
rect 6220 3936 6228 3944
rect 6140 3796 6148 3804
rect 6172 3796 6180 3804
rect 6156 3776 6164 3784
rect 6092 3556 6100 3564
rect 6108 3496 6116 3504
rect 6156 3676 6164 3684
rect 6188 3716 6196 3724
rect 6268 4156 6276 4164
rect 6300 4256 6308 4264
rect 6428 4716 6436 4724
rect 6364 4696 6372 4704
rect 6540 4836 6548 4844
rect 6476 4716 6484 4724
rect 6588 4716 6596 4724
rect 6396 4656 6404 4664
rect 6364 4536 6372 4544
rect 6572 4696 6580 4704
rect 7100 5296 7108 5304
rect 7164 5296 7172 5304
rect 7196 5296 7204 5304
rect 7276 5296 7284 5304
rect 7084 5236 7092 5244
rect 7180 5136 7188 5144
rect 7116 5116 7124 5124
rect 7148 5076 7156 5084
rect 7276 5216 7284 5224
rect 7228 5116 7236 5124
rect 7308 5096 7316 5104
rect 7196 5076 7204 5084
rect 7212 5076 7220 5084
rect 7260 5076 7268 5084
rect 7292 5076 7300 5084
rect 7100 5036 7108 5044
rect 6732 4916 6740 4924
rect 6828 4916 6836 4924
rect 6972 4916 6980 4924
rect 6764 4836 6772 4844
rect 6796 4796 6804 4804
rect 6860 4896 6868 4904
rect 6828 4776 6836 4784
rect 6860 4776 6868 4784
rect 6972 4776 6980 4784
rect 6700 4756 6708 4764
rect 6652 4736 6660 4744
rect 6476 4676 6484 4684
rect 6508 4676 6516 4684
rect 6556 4676 6564 4684
rect 6620 4676 6628 4684
rect 6444 4616 6452 4624
rect 6476 4616 6484 4624
rect 6444 4536 6452 4544
rect 6332 4476 6340 4484
rect 6412 4516 6420 4524
rect 6364 4456 6372 4464
rect 6540 4656 6548 4664
rect 6588 4616 6596 4624
rect 6540 4516 6548 4524
rect 6572 4516 6580 4524
rect 6636 4496 6644 4504
rect 6524 4456 6532 4464
rect 6620 4456 6628 4464
rect 6508 4416 6516 4424
rect 6364 4336 6372 4344
rect 6492 4336 6500 4344
rect 6556 4336 6564 4344
rect 6492 4302 6500 4304
rect 6492 4296 6500 4302
rect 6588 4316 6596 4324
rect 6636 4316 6644 4324
rect 6588 4296 6596 4304
rect 6812 4696 6820 4704
rect 6748 4676 6756 4684
rect 6700 4656 6708 4664
rect 6668 4636 6676 4644
rect 6748 4616 6756 4624
rect 6780 4616 6788 4624
rect 6844 4676 6852 4684
rect 6892 4696 6900 4704
rect 6940 4696 6948 4704
rect 6924 4616 6932 4624
rect 7020 4596 7028 4604
rect 6700 4556 6708 4564
rect 6956 4536 6964 4544
rect 6668 4516 6676 4524
rect 6748 4516 6756 4524
rect 6780 4516 6788 4524
rect 6828 4516 6836 4524
rect 6892 4516 6900 4524
rect 6940 4516 6948 4524
rect 6684 4476 6692 4484
rect 6716 4316 6724 4324
rect 6748 4316 6756 4324
rect 6796 4316 6804 4324
rect 6780 4296 6788 4304
rect 6332 4276 6340 4284
rect 6492 4276 6500 4284
rect 6620 4276 6628 4284
rect 6652 4276 6660 4284
rect 6300 4196 6308 4204
rect 6284 4136 6292 4144
rect 6316 4136 6324 4144
rect 6252 4056 6260 4064
rect 6268 4016 6276 4024
rect 6252 3996 6260 4004
rect 6268 3956 6276 3964
rect 6252 3916 6260 3924
rect 6348 4216 6356 4224
rect 6444 4216 6452 4224
rect 6348 4176 6356 4184
rect 6364 4176 6372 4184
rect 6300 4076 6308 4084
rect 6316 4016 6324 4024
rect 6284 3916 6292 3924
rect 6268 3876 6276 3884
rect 6236 3856 6244 3864
rect 6284 3856 6292 3864
rect 6300 3856 6308 3864
rect 6252 3776 6260 3784
rect 6252 3756 6260 3764
rect 6220 3656 6228 3664
rect 6188 3636 6196 3644
rect 6204 3636 6212 3644
rect 6108 3456 6116 3464
rect 6124 3456 6132 3464
rect 6092 3376 6100 3384
rect 6044 3236 6052 3244
rect 5996 3216 6004 3224
rect 5916 3102 5924 3104
rect 5916 3096 5924 3102
rect 5852 3036 5860 3044
rect 5788 3016 5796 3024
rect 5868 3016 5876 3024
rect 5923 3006 5931 3014
rect 5933 3006 5941 3014
rect 5943 3006 5951 3014
rect 5953 3006 5961 3014
rect 5963 3006 5971 3014
rect 5973 3006 5981 3014
rect 5900 2996 5908 3004
rect 5820 2936 5828 2944
rect 5820 2896 5828 2904
rect 5820 2796 5828 2804
rect 5788 2756 5796 2764
rect 5804 2756 5812 2764
rect 5772 2736 5780 2744
rect 5772 2716 5780 2724
rect 5788 2716 5796 2724
rect 5756 2696 5764 2704
rect 5740 2596 5748 2604
rect 5692 2556 5700 2564
rect 5612 2376 5620 2384
rect 5692 2336 5700 2344
rect 5612 2316 5620 2324
rect 5660 2316 5668 2324
rect 5676 2276 5684 2284
rect 5820 2656 5828 2664
rect 5820 2636 5828 2644
rect 5788 2616 5796 2624
rect 5820 2616 5828 2624
rect 5804 2596 5812 2604
rect 5772 2476 5780 2484
rect 5772 2456 5780 2464
rect 5804 2456 5812 2464
rect 5772 2416 5780 2424
rect 5708 2276 5716 2284
rect 5804 2336 5812 2344
rect 5788 2316 5796 2324
rect 5788 2296 5796 2304
rect 5804 2296 5812 2304
rect 5740 2276 5748 2284
rect 5756 2276 5764 2284
rect 5692 2256 5700 2264
rect 5724 2256 5732 2264
rect 5772 2256 5780 2264
rect 5740 2216 5748 2224
rect 5676 2196 5684 2204
rect 5628 2176 5636 2184
rect 5644 2176 5652 2184
rect 5660 2156 5668 2164
rect 5612 2136 5620 2144
rect 5596 2056 5604 2064
rect 5548 1956 5556 1964
rect 5532 1916 5540 1924
rect 5516 1896 5524 1904
rect 5548 1896 5556 1904
rect 5468 1876 5476 1884
rect 5452 1856 5460 1864
rect 5484 1736 5492 1744
rect 5452 1716 5460 1724
rect 5564 1876 5572 1884
rect 5532 1756 5540 1764
rect 5548 1756 5556 1764
rect 5516 1716 5524 1724
rect 5484 1656 5492 1664
rect 5500 1656 5508 1664
rect 5468 1636 5476 1644
rect 5580 1856 5588 1864
rect 5756 2176 5764 2184
rect 5644 2116 5652 2124
rect 5676 2116 5684 2124
rect 5660 2016 5668 2024
rect 5644 1936 5652 1944
rect 5772 2156 5780 2164
rect 5772 2076 5780 2084
rect 5740 1996 5748 2004
rect 5708 1956 5716 1964
rect 5676 1936 5684 1944
rect 5740 1916 5748 1924
rect 5628 1876 5636 1884
rect 5660 1796 5668 1804
rect 5596 1776 5604 1784
rect 5644 1776 5652 1784
rect 5580 1756 5588 1764
rect 5932 2896 5940 2904
rect 5980 2896 5988 2904
rect 5884 2876 5892 2884
rect 5932 2796 5940 2804
rect 5900 2736 5908 2744
rect 6076 3256 6084 3264
rect 6076 3096 6084 3104
rect 6012 2796 6020 2804
rect 6028 2756 6036 2764
rect 5996 2696 6004 2704
rect 5868 2676 5876 2684
rect 5868 2656 5876 2664
rect 5852 2636 5860 2644
rect 5923 2606 5931 2614
rect 5933 2606 5941 2614
rect 5943 2606 5951 2614
rect 5953 2606 5961 2614
rect 5963 2606 5971 2614
rect 5973 2606 5981 2614
rect 5852 2536 5860 2544
rect 5900 2516 5908 2524
rect 5868 2436 5876 2444
rect 5836 2416 5844 2424
rect 5884 2376 5892 2384
rect 5836 2336 5844 2344
rect 5820 2256 5828 2264
rect 5868 2216 5876 2224
rect 5836 2196 5844 2204
rect 5868 2136 5876 2144
rect 5884 2096 5892 2104
rect 5980 2496 5988 2504
rect 5916 2276 5924 2284
rect 5923 2206 5931 2214
rect 5933 2206 5941 2214
rect 5943 2206 5951 2214
rect 5953 2206 5961 2214
rect 5963 2206 5971 2214
rect 5973 2206 5981 2214
rect 5964 2176 5972 2184
rect 5932 2136 5940 2144
rect 5916 2116 5924 2124
rect 5900 2076 5908 2084
rect 5788 2056 5796 2064
rect 5788 1976 5796 1984
rect 5932 1956 5940 1964
rect 5836 1936 5844 1944
rect 5852 1936 5860 1944
rect 5788 1896 5796 1904
rect 5756 1856 5764 1864
rect 5724 1836 5732 1844
rect 5756 1836 5764 1844
rect 5884 1916 5892 1924
rect 5916 1896 5924 1904
rect 5756 1816 5764 1824
rect 5772 1816 5780 1824
rect 5708 1756 5716 1764
rect 5740 1756 5748 1764
rect 5628 1696 5636 1704
rect 5772 1736 5780 1744
rect 5868 1816 5876 1824
rect 5852 1776 5860 1784
rect 5820 1756 5828 1764
rect 5836 1736 5844 1744
rect 5980 2116 5988 2124
rect 5964 1856 5972 1864
rect 5980 1856 5988 1864
rect 5923 1806 5931 1814
rect 5933 1806 5941 1814
rect 5943 1806 5951 1814
rect 5953 1806 5961 1814
rect 5963 1806 5971 1814
rect 5973 1806 5981 1814
rect 5900 1776 5908 1784
rect 5900 1756 5908 1764
rect 5884 1736 5892 1744
rect 5676 1696 5684 1704
rect 5692 1696 5700 1704
rect 5692 1656 5700 1664
rect 5516 1596 5524 1604
rect 5564 1636 5572 1644
rect 5644 1636 5652 1644
rect 5820 1656 5828 1664
rect 5804 1616 5812 1624
rect 5596 1516 5604 1524
rect 5468 1496 5476 1504
rect 5532 1496 5540 1504
rect 5564 1476 5572 1484
rect 5436 1436 5444 1444
rect 5420 1416 5428 1424
rect 5532 1436 5540 1444
rect 5500 1416 5508 1424
rect 5452 1396 5460 1404
rect 5580 1416 5588 1424
rect 5532 1396 5540 1404
rect 5692 1476 5700 1484
rect 5692 1416 5700 1424
rect 5644 1356 5652 1364
rect 5724 1396 5732 1404
rect 5708 1376 5716 1384
rect 5660 1316 5668 1324
rect 5676 1316 5684 1324
rect 5452 1176 5460 1184
rect 5404 1116 5412 1124
rect 5532 1196 5540 1204
rect 5692 1296 5700 1304
rect 5644 1236 5652 1244
rect 5660 1236 5668 1244
rect 5644 1196 5652 1204
rect 5516 1176 5524 1184
rect 5564 1176 5572 1184
rect 5596 1176 5604 1184
rect 5468 1156 5476 1164
rect 5484 1116 5492 1124
rect 5500 1116 5508 1124
rect 5340 1096 5348 1104
rect 5356 1096 5364 1104
rect 5388 1096 5396 1104
rect 5324 1076 5332 1084
rect 5436 1076 5444 1084
rect 5420 1056 5428 1064
rect 5372 1036 5380 1044
rect 5404 1036 5412 1044
rect 5388 996 5396 1004
rect 5308 956 5316 964
rect 5276 936 5284 944
rect 5452 956 5460 964
rect 5468 956 5476 964
rect 5580 1116 5588 1124
rect 5516 1076 5524 1084
rect 5532 1056 5540 1064
rect 5516 1016 5524 1024
rect 5500 956 5508 964
rect 5452 936 5460 944
rect 5484 936 5492 944
rect 5548 976 5556 984
rect 5532 956 5540 964
rect 5676 1176 5684 1184
rect 5660 1096 5668 1104
rect 5708 1256 5716 1264
rect 5868 1596 5876 1604
rect 6028 2536 6036 2544
rect 6012 2516 6020 2524
rect 6028 2476 6036 2484
rect 6076 3056 6084 3064
rect 6092 3036 6100 3044
rect 6076 3016 6084 3024
rect 6156 3436 6164 3444
rect 6220 3516 6228 3524
rect 6220 3502 6228 3504
rect 6220 3496 6228 3502
rect 6220 3456 6228 3464
rect 6188 3356 6196 3364
rect 6124 3336 6132 3344
rect 6156 3316 6164 3324
rect 6188 3256 6196 3264
rect 6124 3036 6132 3044
rect 6092 2956 6100 2964
rect 6108 2836 6116 2844
rect 6108 2736 6116 2744
rect 6172 3076 6180 3084
rect 6204 3056 6212 3064
rect 6188 2976 6196 2984
rect 6156 2876 6164 2884
rect 6140 2856 6148 2864
rect 6140 2696 6148 2704
rect 6412 4136 6420 4144
rect 6428 4056 6436 4064
rect 6476 4096 6484 4104
rect 6460 4036 6468 4044
rect 6396 3996 6404 4004
rect 6380 3936 6388 3944
rect 6364 3916 6372 3924
rect 6316 3716 6324 3724
rect 6300 3676 6308 3684
rect 6348 3776 6356 3784
rect 6380 3756 6388 3764
rect 6412 3936 6420 3944
rect 6444 3916 6452 3924
rect 6412 3816 6420 3824
rect 6476 3996 6484 4004
rect 6524 4256 6532 4264
rect 6508 4196 6516 4204
rect 6572 4196 6580 4204
rect 6540 4116 6548 4124
rect 6508 4076 6516 4084
rect 6508 3936 6516 3944
rect 6556 4096 6564 4104
rect 6588 4076 6596 4084
rect 6572 4016 6580 4024
rect 6652 4256 6660 4264
rect 6652 4076 6660 4084
rect 6620 3976 6628 3984
rect 6572 3936 6580 3944
rect 6508 3916 6516 3924
rect 6540 3916 6548 3924
rect 6892 4316 6900 4324
rect 6812 4276 6820 4284
rect 6844 4276 6852 4284
rect 6956 4276 6964 4284
rect 6716 4236 6724 4244
rect 6828 4196 6836 4204
rect 6812 4156 6820 4164
rect 6748 4136 6756 4144
rect 6700 4096 6708 4104
rect 6796 4096 6804 4104
rect 6780 4076 6788 4084
rect 6668 3976 6676 3984
rect 6684 3956 6692 3964
rect 6748 3936 6756 3944
rect 6492 3896 6500 3904
rect 6652 3896 6660 3904
rect 6492 3876 6500 3884
rect 6492 3856 6500 3864
rect 6396 3736 6404 3744
rect 6476 3736 6484 3744
rect 6620 3876 6628 3884
rect 6540 3856 6548 3864
rect 6556 3816 6564 3824
rect 6812 3916 6820 3924
rect 6828 3916 6836 3924
rect 6780 3896 6788 3904
rect 6668 3876 6676 3884
rect 6700 3856 6708 3864
rect 6620 3836 6628 3844
rect 6636 3836 6644 3844
rect 6572 3796 6580 3804
rect 6428 3696 6436 3704
rect 6348 3676 6356 3684
rect 6332 3656 6340 3664
rect 6492 3596 6500 3604
rect 6348 3556 6356 3564
rect 6396 3556 6404 3564
rect 6364 3536 6372 3544
rect 6412 3496 6420 3504
rect 6252 3416 6260 3424
rect 6316 3396 6324 3404
rect 6380 3356 6388 3364
rect 6348 3316 6356 3324
rect 6236 3116 6244 3124
rect 6476 3416 6484 3424
rect 6444 3396 6452 3404
rect 6412 3336 6420 3344
rect 6460 3336 6468 3344
rect 6444 3256 6452 3264
rect 6588 3716 6596 3724
rect 6540 3696 6548 3704
rect 6732 3836 6740 3844
rect 6716 3776 6724 3784
rect 6652 3736 6660 3744
rect 6668 3716 6676 3724
rect 6620 3696 6628 3704
rect 6652 3696 6660 3704
rect 6716 3716 6724 3724
rect 6764 3696 6772 3704
rect 6604 3676 6612 3684
rect 6700 3676 6708 3684
rect 6828 3896 6836 3904
rect 6940 4236 6948 4244
rect 6924 4216 6932 4224
rect 6908 4176 6916 4184
rect 6924 4176 6932 4184
rect 6972 4176 6980 4184
rect 6876 4116 6884 4124
rect 6940 4096 6948 4104
rect 6940 4076 6948 4084
rect 6924 4036 6932 4044
rect 6892 4016 6900 4024
rect 6860 3936 6868 3944
rect 6892 3876 6900 3884
rect 6844 3756 6852 3764
rect 6844 3736 6852 3744
rect 6796 3716 6804 3724
rect 6812 3716 6820 3724
rect 6796 3656 6804 3664
rect 6716 3616 6724 3624
rect 6780 3616 6788 3624
rect 6828 3616 6836 3624
rect 6636 3536 6644 3544
rect 6684 3536 6692 3544
rect 6540 3516 6548 3524
rect 6652 3516 6660 3524
rect 6604 3496 6612 3504
rect 6748 3496 6756 3504
rect 6876 3696 6884 3704
rect 6876 3556 6884 3564
rect 6860 3516 6868 3524
rect 6492 3376 6500 3384
rect 6540 3336 6548 3344
rect 6572 3316 6580 3324
rect 6652 3316 6660 3324
rect 6476 3276 6484 3284
rect 6492 3256 6500 3264
rect 6588 3236 6596 3244
rect 6668 3236 6676 3244
rect 6460 3156 6468 3164
rect 6572 3176 6580 3184
rect 6476 3116 6484 3124
rect 6524 3116 6532 3124
rect 6572 3116 6580 3124
rect 6268 3096 6276 3104
rect 6332 3096 6340 3104
rect 6396 3096 6404 3104
rect 6524 3096 6532 3104
rect 6300 3076 6308 3084
rect 6316 3056 6324 3064
rect 6460 3076 6468 3084
rect 6364 3036 6372 3044
rect 6364 3016 6372 3024
rect 6300 2996 6308 3004
rect 6332 2996 6340 3004
rect 6380 2956 6388 2964
rect 6412 2956 6420 2964
rect 6348 2916 6356 2924
rect 6460 3036 6468 3044
rect 6476 3036 6484 3044
rect 6204 2896 6212 2904
rect 6204 2716 6212 2724
rect 6124 2676 6132 2684
rect 6060 2616 6068 2624
rect 6140 2616 6148 2624
rect 6124 2596 6132 2604
rect 6124 2556 6132 2564
rect 6108 2536 6116 2544
rect 6092 2476 6100 2484
rect 6140 2456 6148 2464
rect 6044 2376 6052 2384
rect 6060 2376 6068 2384
rect 6076 2376 6084 2384
rect 6060 2256 6068 2264
rect 6060 2216 6068 2224
rect 6028 2156 6036 2164
rect 6060 2076 6068 2084
rect 6044 1996 6052 2004
rect 6028 1976 6036 1984
rect 6012 1916 6020 1924
rect 6044 1896 6052 1904
rect 6108 2316 6116 2324
rect 6092 2296 6100 2304
rect 6172 2676 6180 2684
rect 6188 2676 6196 2684
rect 6156 2316 6164 2324
rect 6140 2196 6148 2204
rect 6124 2136 6132 2144
rect 6092 2116 6100 2124
rect 6092 2036 6100 2044
rect 6076 2016 6084 2024
rect 6140 2116 6148 2124
rect 6124 2036 6132 2044
rect 6108 1996 6116 2004
rect 6092 1976 6100 1984
rect 6092 1936 6100 1944
rect 6124 1936 6132 1944
rect 6076 1916 6084 1924
rect 6108 1856 6116 1864
rect 6076 1816 6084 1824
rect 6092 1796 6100 1804
rect 6076 1776 6084 1784
rect 5900 1596 5908 1604
rect 5900 1556 5908 1564
rect 6060 1736 6068 1744
rect 6060 1716 6068 1724
rect 5996 1656 6004 1664
rect 6044 1636 6052 1644
rect 5996 1616 6004 1624
rect 5996 1536 6004 1544
rect 5900 1516 5908 1524
rect 5916 1516 5924 1524
rect 5980 1516 5988 1524
rect 5804 1476 5812 1484
rect 5852 1476 5860 1484
rect 5772 1376 5780 1384
rect 5788 1376 5796 1384
rect 5772 1356 5780 1364
rect 5788 1316 5796 1324
rect 5740 1196 5748 1204
rect 5724 1176 5732 1184
rect 5788 1156 5796 1164
rect 5724 1136 5732 1144
rect 5708 1116 5716 1124
rect 5772 1116 5780 1124
rect 5708 1096 5716 1104
rect 5692 1076 5700 1084
rect 5724 1056 5732 1064
rect 5676 1016 5684 1024
rect 5580 956 5588 964
rect 5564 936 5572 944
rect 5660 936 5668 944
rect 5500 916 5508 924
rect 5196 796 5204 804
rect 5260 796 5268 804
rect 5036 776 5044 784
rect 5116 776 5124 784
rect 4956 736 4964 744
rect 5340 896 5348 904
rect 5356 836 5364 844
rect 5308 756 5316 764
rect 5324 736 5332 744
rect 4956 696 4964 704
rect 5020 702 5028 704
rect 5020 696 5028 702
rect 4924 676 4932 684
rect 4940 616 4948 624
rect 4924 576 4932 584
rect 4908 556 4916 564
rect 4908 476 4916 484
rect 5084 676 5092 684
rect 5164 696 5172 704
rect 5244 696 5252 704
rect 5148 656 5156 664
rect 5260 656 5268 664
rect 5116 616 5124 624
rect 5212 596 5220 604
rect 5388 702 5396 704
rect 5388 696 5396 702
rect 5292 616 5300 624
rect 5372 616 5380 624
rect 5116 556 5124 564
rect 5180 556 5188 564
rect 5212 556 5220 564
rect 5228 556 5236 564
rect 5308 556 5316 564
rect 5484 896 5492 904
rect 5452 796 5460 804
rect 5516 896 5524 904
rect 5756 1076 5764 1084
rect 5612 916 5620 924
rect 5708 916 5716 924
rect 5564 896 5572 904
rect 5548 796 5556 804
rect 5548 756 5556 764
rect 5532 736 5540 744
rect 5500 696 5508 704
rect 5452 676 5460 684
rect 5404 596 5412 604
rect 5468 556 5476 564
rect 5404 536 5412 544
rect 5484 536 5492 544
rect 4956 496 4964 504
rect 4956 476 4964 484
rect 4940 436 4948 444
rect 5052 518 5060 524
rect 5052 516 5060 518
rect 5148 496 5156 504
rect 5116 476 5124 484
rect 5020 456 5028 464
rect 4972 436 4980 444
rect 4940 356 4948 364
rect 4956 356 4964 364
rect 4908 316 4916 324
rect 4876 276 4884 284
rect 4892 276 4900 284
rect 4924 256 4932 264
rect 4796 176 4804 184
rect 4924 236 4932 244
rect 4844 196 4852 204
rect 4860 196 4868 204
rect 4908 176 4916 184
rect 4924 176 4932 184
rect 4828 76 4836 84
rect 4860 76 4868 84
rect 4892 36 4900 44
rect 5068 276 5076 284
rect 4972 256 4980 264
rect 4956 236 4964 244
rect 4988 236 4996 244
rect 5196 516 5204 524
rect 5212 496 5220 504
rect 5212 456 5220 464
rect 5180 336 5188 344
rect 5148 316 5156 324
rect 5164 296 5172 304
rect 5132 276 5140 284
rect 5148 236 5156 244
rect 5052 156 5060 164
rect 5004 136 5012 144
rect 5036 116 5044 124
rect 5068 96 5076 104
rect 5116 116 5124 124
rect 5196 216 5204 224
rect 5260 516 5268 524
rect 5324 516 5332 524
rect 5388 516 5396 524
rect 5276 356 5284 364
rect 5244 336 5252 344
rect 5228 236 5236 244
rect 5468 516 5476 524
rect 5436 476 5444 484
rect 5436 316 5444 324
rect 5340 256 5348 264
rect 5276 216 5284 224
rect 5308 216 5316 224
rect 5628 796 5636 804
rect 5644 676 5652 684
rect 5580 616 5588 624
rect 5740 656 5748 664
rect 5788 676 5796 684
rect 5772 636 5780 644
rect 5676 616 5684 624
rect 5708 616 5716 624
rect 5740 616 5748 624
rect 5772 616 5780 624
rect 5372 256 5380 264
rect 5436 256 5444 264
rect 5484 256 5492 264
rect 5468 196 5476 204
rect 5356 176 5364 184
rect 5276 136 5284 144
rect 5548 136 5556 144
rect 5788 556 5796 564
rect 5868 1436 5876 1444
rect 5884 1396 5892 1404
rect 5923 1406 5931 1414
rect 5933 1406 5941 1414
rect 5943 1406 5951 1414
rect 5953 1406 5961 1414
rect 5963 1406 5971 1414
rect 5973 1406 5981 1414
rect 5948 1356 5956 1364
rect 5884 1196 5892 1204
rect 5820 1176 5828 1184
rect 5868 1156 5876 1164
rect 5836 1096 5844 1104
rect 5852 1076 5860 1084
rect 5836 1036 5844 1044
rect 5820 756 5828 764
rect 5884 1096 5892 1104
rect 5916 1316 5924 1324
rect 5980 1176 5988 1184
rect 5916 1116 5924 1124
rect 5923 1006 5931 1014
rect 5933 1006 5941 1014
rect 5943 1006 5951 1014
rect 5953 1006 5961 1014
rect 5963 1006 5971 1014
rect 5973 1006 5981 1014
rect 6188 2276 6196 2284
rect 6172 2256 6180 2264
rect 6172 2196 6180 2204
rect 6316 2896 6324 2904
rect 6364 2896 6372 2904
rect 6380 2896 6388 2904
rect 6252 2876 6260 2884
rect 6300 2776 6308 2784
rect 6268 2696 6276 2704
rect 6252 2636 6260 2644
rect 6252 2476 6260 2484
rect 6364 2876 6372 2884
rect 6332 2776 6340 2784
rect 6316 2676 6324 2684
rect 6316 2636 6324 2644
rect 6396 2876 6404 2884
rect 6396 2736 6404 2744
rect 6396 2656 6404 2664
rect 6364 2636 6372 2644
rect 6428 2896 6436 2904
rect 6460 2876 6468 2884
rect 6460 2696 6468 2704
rect 6428 2676 6436 2684
rect 6460 2676 6468 2684
rect 6604 3096 6612 3104
rect 6556 3076 6564 3084
rect 6540 2996 6548 3004
rect 6636 3076 6644 3084
rect 6588 3056 6596 3064
rect 6572 3016 6580 3024
rect 6556 2916 6564 2924
rect 6508 2856 6516 2864
rect 6524 2676 6532 2684
rect 6492 2656 6500 2664
rect 6412 2616 6420 2624
rect 6300 2556 6308 2564
rect 6364 2536 6372 2544
rect 6508 2616 6516 2624
rect 6556 2656 6564 2664
rect 6444 2576 6452 2584
rect 6364 2516 6372 2524
rect 6380 2516 6388 2524
rect 6316 2376 6324 2384
rect 6284 2316 6292 2324
rect 6300 2316 6308 2324
rect 6220 2296 6228 2304
rect 6236 2296 6244 2304
rect 6284 2296 6292 2304
rect 6236 2216 6244 2224
rect 6268 2176 6276 2184
rect 6204 2156 6212 2164
rect 6252 2136 6260 2144
rect 6172 2096 6180 2104
rect 6172 2076 6180 2084
rect 6156 1956 6164 1964
rect 6140 1916 6148 1924
rect 6140 1896 6148 1904
rect 6156 1856 6164 1864
rect 6236 1996 6244 2004
rect 6188 1896 6196 1904
rect 6172 1836 6180 1844
rect 6124 1756 6132 1764
rect 6172 1736 6180 1744
rect 6140 1636 6148 1644
rect 6076 1616 6084 1624
rect 6108 1596 6116 1604
rect 6060 1556 6068 1564
rect 6092 1556 6100 1564
rect 6028 1536 6036 1544
rect 6044 1516 6052 1524
rect 6140 1516 6148 1524
rect 6092 1496 6100 1504
rect 6124 1496 6132 1504
rect 6140 1436 6148 1444
rect 6076 1416 6084 1424
rect 6108 1396 6116 1404
rect 6060 1356 6068 1364
rect 6012 1336 6020 1344
rect 6044 1336 6052 1344
rect 6028 1296 6036 1304
rect 6012 1216 6020 1224
rect 6060 1276 6068 1284
rect 6044 1256 6052 1264
rect 6108 1296 6116 1304
rect 6108 1276 6116 1284
rect 6092 1216 6100 1224
rect 6076 1196 6084 1204
rect 6060 1176 6068 1184
rect 6028 1036 6036 1044
rect 5900 916 5908 924
rect 5900 896 5908 904
rect 5836 676 5844 684
rect 5868 656 5876 664
rect 5884 636 5892 644
rect 5868 576 5876 584
rect 5596 516 5604 524
rect 5708 516 5716 524
rect 5788 516 5796 524
rect 5820 516 5828 524
rect 5612 476 5620 484
rect 5596 316 5604 324
rect 5804 496 5812 504
rect 5820 476 5828 484
rect 5788 336 5796 344
rect 5740 316 5748 324
rect 5788 316 5796 324
rect 5644 296 5652 304
rect 5660 296 5668 304
rect 5836 316 5844 324
rect 5980 856 5988 864
rect 5996 796 6004 804
rect 6012 796 6020 804
rect 5932 676 5940 684
rect 6012 756 6020 764
rect 5996 656 6004 664
rect 5923 606 5931 614
rect 5933 606 5941 614
rect 5943 606 5951 614
rect 5953 606 5961 614
rect 5963 606 5971 614
rect 5973 606 5981 614
rect 5900 596 5908 604
rect 6060 1076 6068 1084
rect 6092 1176 6100 1184
rect 6092 1076 6100 1084
rect 6204 1856 6212 1864
rect 6220 1856 6228 1864
rect 6268 2116 6276 2124
rect 6492 2536 6500 2544
rect 6508 2536 6516 2544
rect 6540 2576 6548 2584
rect 6556 2536 6564 2544
rect 6428 2496 6436 2504
rect 6444 2496 6452 2504
rect 6492 2496 6500 2504
rect 6444 2456 6452 2464
rect 6412 2376 6420 2384
rect 6380 2316 6388 2324
rect 6332 2296 6340 2304
rect 6380 2276 6388 2284
rect 6364 2256 6372 2264
rect 6364 2176 6372 2184
rect 6412 2176 6420 2184
rect 6332 2076 6340 2084
rect 6300 2016 6308 2024
rect 6332 2016 6340 2024
rect 6268 1896 6276 1904
rect 6284 1896 6292 1904
rect 6284 1856 6292 1864
rect 6284 1796 6292 1804
rect 6204 1756 6212 1764
rect 6220 1756 6228 1764
rect 6252 1736 6260 1744
rect 6220 1716 6228 1724
rect 6268 1716 6276 1724
rect 6700 3436 6708 3444
rect 6812 3476 6820 3484
rect 6764 3376 6772 3384
rect 6844 3456 6852 3464
rect 6844 3376 6852 3384
rect 6796 3296 6804 3304
rect 6684 3136 6692 3144
rect 6652 3036 6660 3044
rect 6620 2976 6628 2984
rect 6620 2936 6628 2944
rect 6604 2856 6612 2864
rect 6604 2716 6612 2724
rect 6604 2696 6612 2704
rect 6652 2916 6660 2924
rect 6668 2876 6676 2884
rect 6700 3116 6708 3124
rect 6700 2996 6708 3004
rect 6748 3116 6756 3124
rect 6700 2896 6708 2904
rect 6732 2896 6740 2904
rect 6684 2656 6692 2664
rect 6636 2636 6644 2644
rect 6620 2596 6628 2604
rect 6588 2576 6596 2584
rect 6684 2556 6692 2564
rect 6652 2496 6660 2504
rect 6540 2436 6548 2444
rect 6476 2416 6484 2424
rect 6460 2396 6468 2404
rect 6444 2296 6452 2304
rect 6460 2296 6468 2304
rect 6444 2116 6452 2124
rect 6460 2116 6468 2124
rect 6428 1996 6436 2004
rect 6540 2336 6548 2344
rect 6492 2316 6500 2324
rect 6508 2236 6516 2244
rect 6524 2236 6532 2244
rect 6716 2736 6724 2744
rect 6828 3256 6836 3264
rect 6908 3776 6916 3784
rect 6940 3856 6948 3864
rect 7180 4976 7188 4984
rect 7100 4956 7108 4964
rect 7052 4936 7060 4944
rect 7084 4616 7092 4624
rect 7068 4596 7076 4604
rect 7132 4896 7140 4904
rect 7148 4736 7156 4744
rect 7132 4696 7140 4704
rect 7164 4636 7172 4644
rect 7164 4596 7172 4604
rect 7100 4536 7108 4544
rect 7132 4516 7140 4524
rect 7052 4296 7060 4304
rect 7148 4496 7156 4504
rect 7340 5036 7348 5044
rect 7212 4956 7220 4964
rect 7292 4916 7300 4924
rect 7228 4696 7236 4704
rect 7180 4456 7188 4464
rect 7180 4316 7188 4324
rect 7180 4296 7188 4304
rect 7132 4276 7140 4284
rect 7148 4276 7156 4284
rect 7180 4276 7188 4284
rect 7052 4136 7060 4144
rect 7084 4116 7092 4124
rect 7036 4096 7044 4104
rect 6972 3916 6980 3924
rect 6956 3836 6964 3844
rect 6940 3816 6948 3824
rect 6924 3736 6932 3744
rect 6924 3656 6932 3664
rect 6908 3636 6916 3644
rect 6892 3536 6900 3544
rect 6924 3556 6932 3564
rect 6924 3536 6932 3544
rect 6892 3476 6900 3484
rect 6876 3456 6884 3464
rect 6908 3436 6916 3444
rect 6908 3316 6916 3324
rect 6876 3136 6884 3144
rect 6812 3056 6820 3064
rect 6812 3016 6820 3024
rect 6860 3076 6868 3084
rect 6876 3076 6884 3084
rect 6844 2996 6852 3004
rect 6780 2976 6788 2984
rect 6764 2836 6772 2844
rect 6748 2636 6756 2644
rect 6796 2716 6804 2724
rect 6908 3036 6916 3044
rect 6892 2956 6900 2964
rect 6908 2876 6916 2884
rect 6924 2776 6932 2784
rect 6892 2736 6900 2744
rect 6924 2736 6932 2744
rect 6876 2696 6884 2704
rect 6892 2676 6900 2684
rect 6844 2656 6852 2664
rect 6876 2616 6884 2624
rect 6764 2596 6772 2604
rect 6860 2596 6868 2604
rect 6748 2576 6756 2584
rect 6732 2516 6740 2524
rect 6700 2416 6708 2424
rect 6620 2396 6628 2404
rect 6700 2396 6708 2404
rect 6556 2316 6564 2324
rect 6572 2316 6580 2324
rect 6700 2376 6708 2384
rect 6636 2296 6644 2304
rect 6652 2296 6660 2304
rect 6684 2296 6692 2304
rect 6556 2276 6564 2284
rect 6604 2236 6612 2244
rect 6588 2216 6596 2224
rect 6668 2276 6676 2284
rect 6652 2256 6660 2264
rect 6716 2236 6724 2244
rect 6620 2196 6628 2204
rect 6684 2196 6692 2204
rect 6556 2176 6564 2184
rect 6508 2116 6516 2124
rect 6492 1936 6500 1944
rect 6492 1916 6500 1924
rect 6348 1876 6356 1884
rect 6396 1876 6404 1884
rect 6412 1876 6420 1884
rect 6332 1796 6340 1804
rect 6476 1876 6484 1884
rect 6508 1880 6516 1884
rect 6508 1876 6516 1880
rect 6540 2036 6548 2044
rect 6540 1996 6548 2004
rect 6636 2156 6644 2164
rect 6588 2136 6596 2144
rect 6732 2196 6740 2204
rect 6620 2116 6628 2124
rect 6572 2096 6580 2104
rect 6716 2096 6724 2104
rect 6684 2076 6692 2084
rect 6620 1976 6628 1984
rect 6668 1976 6676 1984
rect 6604 1936 6612 1944
rect 6572 1876 6580 1884
rect 6428 1836 6436 1844
rect 6460 1836 6468 1844
rect 6380 1816 6388 1824
rect 6428 1816 6436 1824
rect 6316 1756 6324 1764
rect 6364 1756 6372 1764
rect 6300 1736 6308 1744
rect 6364 1736 6372 1744
rect 6412 1756 6420 1764
rect 6508 1856 6516 1864
rect 6524 1856 6532 1864
rect 6492 1756 6500 1764
rect 6556 1816 6564 1824
rect 6588 1796 6596 1804
rect 6540 1756 6548 1764
rect 6556 1736 6564 1744
rect 6300 1716 6308 1724
rect 6476 1716 6484 1724
rect 6732 1916 6740 1924
rect 6652 1876 6660 1884
rect 6876 2576 6884 2584
rect 6812 2516 6820 2524
rect 6812 2496 6820 2504
rect 6844 2496 6852 2504
rect 6876 2456 6884 2464
rect 6812 2296 6820 2304
rect 6796 2256 6804 2264
rect 6780 2136 6788 2144
rect 6860 2376 6868 2384
rect 6860 2316 6868 2324
rect 6844 2236 6852 2244
rect 6844 2196 6852 2204
rect 6828 2116 6836 2124
rect 6764 2096 6772 2104
rect 6780 2056 6788 2064
rect 6668 1816 6676 1824
rect 6748 1816 6756 1824
rect 6652 1796 6660 1804
rect 6636 1756 6644 1764
rect 6604 1736 6612 1744
rect 6620 1736 6628 1744
rect 6764 1776 6772 1784
rect 6748 1736 6756 1744
rect 6652 1716 6660 1724
rect 6284 1676 6292 1684
rect 6300 1676 6308 1684
rect 6204 1576 6212 1584
rect 6236 1576 6244 1584
rect 6188 1556 6196 1564
rect 6220 1556 6228 1564
rect 6188 1476 6196 1484
rect 6204 1456 6212 1464
rect 6172 1436 6180 1444
rect 6204 1416 6212 1424
rect 6284 1516 6292 1524
rect 6316 1656 6324 1664
rect 6444 1696 6452 1704
rect 6348 1536 6356 1544
rect 6396 1516 6404 1524
rect 6332 1496 6340 1504
rect 6588 1696 6596 1704
rect 6444 1636 6452 1644
rect 6492 1636 6500 1644
rect 6476 1556 6484 1564
rect 6572 1616 6580 1624
rect 6588 1616 6596 1624
rect 6620 1596 6628 1604
rect 6508 1576 6516 1584
rect 6524 1576 6532 1584
rect 6460 1496 6468 1504
rect 6364 1476 6372 1484
rect 6412 1476 6420 1484
rect 6444 1476 6452 1484
rect 6252 1456 6260 1464
rect 6268 1456 6276 1464
rect 6316 1456 6324 1464
rect 6236 1416 6244 1424
rect 6348 1416 6356 1424
rect 6172 1356 6180 1364
rect 6332 1376 6340 1384
rect 6348 1376 6356 1384
rect 6156 1296 6164 1304
rect 6492 1476 6500 1484
rect 6380 1456 6388 1464
rect 6460 1456 6468 1464
rect 6396 1376 6404 1384
rect 6412 1376 6420 1384
rect 6460 1376 6468 1384
rect 6476 1376 6484 1384
rect 6492 1376 6500 1384
rect 6396 1356 6404 1364
rect 6428 1356 6436 1364
rect 6220 1236 6228 1244
rect 6172 1216 6180 1224
rect 6204 1196 6212 1204
rect 6140 1156 6148 1164
rect 6156 1156 6164 1164
rect 6188 1136 6196 1144
rect 6172 1096 6180 1104
rect 6140 1076 6148 1084
rect 6220 1096 6228 1104
rect 6284 1296 6292 1304
rect 6252 1216 6260 1224
rect 6268 1196 6276 1204
rect 6108 1036 6116 1044
rect 6140 1036 6148 1044
rect 6044 1016 6052 1024
rect 6076 1016 6084 1024
rect 6140 1016 6148 1024
rect 6156 1016 6164 1024
rect 6044 996 6052 1004
rect 6124 996 6132 1004
rect 6124 936 6132 944
rect 6236 1056 6244 1064
rect 6188 1016 6196 1024
rect 6204 1016 6212 1024
rect 6188 956 6196 964
rect 6076 916 6084 924
rect 6156 916 6164 924
rect 6076 876 6084 884
rect 6060 796 6068 804
rect 5948 556 5956 564
rect 6028 556 6036 564
rect 6012 496 6020 504
rect 6108 756 6116 764
rect 6252 996 6260 1004
rect 6236 976 6244 984
rect 6268 956 6276 964
rect 6220 816 6228 824
rect 6236 796 6244 804
rect 6252 776 6260 784
rect 6140 716 6148 724
rect 6172 716 6180 724
rect 6188 696 6196 704
rect 6204 696 6212 704
rect 6124 676 6132 684
rect 6156 576 6164 584
rect 6140 556 6148 564
rect 6268 736 6276 744
rect 6364 1296 6372 1304
rect 6316 1276 6324 1284
rect 6396 1276 6404 1284
rect 6492 1336 6500 1344
rect 6460 1256 6468 1264
rect 6460 1236 6468 1244
rect 6460 1196 6468 1204
rect 6428 1176 6436 1184
rect 6380 1136 6388 1144
rect 6364 1116 6372 1124
rect 6300 1056 6308 1064
rect 6332 1016 6340 1024
rect 6300 816 6308 824
rect 6284 716 6292 724
rect 6332 856 6340 864
rect 6252 656 6260 664
rect 6060 376 6068 384
rect 6012 336 6020 344
rect 5884 316 5892 324
rect 5996 316 6004 324
rect 5660 216 5668 224
rect 5644 196 5652 204
rect 5660 176 5668 184
rect 5788 256 5796 264
rect 5740 236 5748 244
rect 5708 196 5716 204
rect 5820 176 5828 184
rect 5708 156 5716 164
rect 5884 256 5892 264
rect 5996 256 6004 264
rect 5923 206 5931 214
rect 5933 206 5941 214
rect 5943 206 5951 214
rect 5953 206 5961 214
rect 5963 206 5971 214
rect 5973 206 5981 214
rect 5868 196 5876 204
rect 5900 196 5908 204
rect 5692 136 5700 144
rect 5724 136 5732 144
rect 5836 136 5844 144
rect 6204 376 6212 384
rect 6364 836 6372 844
rect 6492 1116 6500 1124
rect 6428 1056 6436 1064
rect 6396 976 6404 984
rect 6556 1496 6564 1504
rect 6540 1436 6548 1444
rect 6588 1436 6596 1444
rect 6524 1276 6532 1284
rect 6668 1696 6676 1704
rect 6700 1716 6708 1724
rect 6732 1716 6740 1724
rect 6684 1656 6692 1664
rect 6700 1616 6708 1624
rect 6764 1576 6772 1584
rect 6652 1556 6660 1564
rect 6716 1556 6724 1564
rect 6636 1476 6644 1484
rect 6636 1396 6644 1404
rect 6684 1436 6692 1444
rect 6668 1396 6676 1404
rect 6652 1356 6660 1364
rect 6572 1316 6580 1324
rect 6588 1296 6596 1304
rect 6620 1296 6628 1304
rect 6572 1236 6580 1244
rect 6556 1216 6564 1224
rect 6572 1196 6580 1204
rect 6556 1156 6564 1164
rect 6540 1116 6548 1124
rect 6524 1096 6532 1104
rect 6572 1136 6580 1144
rect 6460 1016 6468 1024
rect 6508 1016 6516 1024
rect 6428 956 6436 964
rect 6412 896 6420 904
rect 6412 716 6420 724
rect 6364 636 6372 644
rect 6332 576 6340 584
rect 6348 576 6356 584
rect 6284 518 6292 524
rect 6284 516 6292 518
rect 6444 856 6452 864
rect 6444 616 6452 624
rect 6444 576 6452 584
rect 6508 976 6516 984
rect 6524 936 6532 944
rect 6476 916 6484 924
rect 6508 876 6516 884
rect 6684 1356 6692 1364
rect 6604 976 6612 984
rect 6620 956 6628 964
rect 6540 916 6548 924
rect 6620 916 6628 924
rect 6572 856 6580 864
rect 6476 716 6484 724
rect 6604 776 6612 784
rect 6556 696 6564 704
rect 6604 696 6612 704
rect 6476 676 6484 684
rect 6540 676 6548 684
rect 6588 676 6596 684
rect 6492 656 6500 664
rect 6540 636 6548 644
rect 6556 636 6564 644
rect 6428 536 6436 544
rect 6460 536 6468 544
rect 6380 516 6388 524
rect 6380 496 6388 504
rect 6428 496 6436 504
rect 6396 356 6404 364
rect 6364 336 6372 344
rect 6284 316 6292 324
rect 6332 316 6340 324
rect 6348 316 6356 324
rect 6092 296 6100 304
rect 6140 296 6148 304
rect 6220 296 6228 304
rect 6268 256 6276 264
rect 6220 216 6228 224
rect 6092 176 6100 184
rect 6012 136 6020 144
rect 6060 136 6068 144
rect 5180 116 5188 124
rect 5276 116 5284 124
rect 5340 118 5348 124
rect 5340 116 5348 118
rect 5404 116 5412 124
rect 5580 116 5588 124
rect 5692 116 5700 124
rect 5788 118 5796 124
rect 5788 116 5796 118
rect 5852 116 5860 124
rect 6092 116 6100 124
rect 6284 176 6292 184
rect 6428 316 6436 324
rect 6636 696 6644 704
rect 6524 516 6532 524
rect 6492 496 6500 504
rect 6476 296 6484 304
rect 6476 256 6484 264
rect 6412 216 6420 224
rect 6620 518 6628 524
rect 6620 516 6628 518
rect 6556 496 6564 504
rect 6556 336 6564 344
rect 6572 296 6580 304
rect 6540 236 6548 244
rect 6684 1096 6692 1104
rect 6764 1496 6772 1504
rect 6732 1476 6740 1484
rect 6732 1456 6740 1464
rect 6812 2036 6820 2044
rect 6844 1976 6852 1984
rect 6924 2616 6932 2624
rect 6908 2496 6916 2504
rect 6892 2296 6900 2304
rect 7084 4096 7092 4104
rect 7164 4076 7172 4084
rect 7132 4056 7140 4064
rect 7260 4116 7268 4124
rect 7196 4016 7204 4024
rect 7212 4016 7220 4024
rect 7148 3916 7156 3924
rect 7180 3916 7188 3924
rect 7100 3896 7108 3904
rect 7148 3896 7156 3904
rect 7196 3896 7204 3904
rect 7020 3876 7028 3884
rect 7052 3856 7060 3864
rect 7084 3856 7092 3864
rect 7036 3816 7044 3824
rect 6988 3796 6996 3804
rect 7004 3756 7012 3764
rect 6972 3696 6980 3704
rect 7020 3656 7028 3664
rect 6988 3616 6996 3624
rect 7004 3616 7012 3624
rect 7020 3556 7028 3564
rect 7020 3516 7028 3524
rect 7084 3796 7092 3804
rect 7068 3776 7076 3784
rect 7052 3736 7060 3744
rect 7068 3656 7076 3664
rect 7052 3596 7060 3604
rect 7004 3456 7012 3464
rect 7036 3456 7044 3464
rect 6956 3296 6964 3304
rect 6972 3256 6980 3264
rect 6956 3176 6964 3184
rect 6956 3136 6964 3144
rect 6988 3236 6996 3244
rect 6988 3056 6996 3064
rect 6972 2976 6980 2984
rect 7036 3436 7044 3444
rect 7052 3316 7060 3324
rect 7036 3256 7044 3264
rect 7020 3116 7028 3124
rect 7036 3096 7044 3104
rect 7004 2976 7012 2984
rect 7020 2956 7028 2964
rect 6988 2936 6996 2944
rect 7004 2916 7012 2924
rect 7004 2736 7012 2744
rect 6972 2716 6980 2724
rect 6972 2696 6980 2704
rect 7020 2636 7028 2644
rect 6988 2596 6996 2604
rect 7004 2596 7012 2604
rect 6988 2576 6996 2584
rect 6956 2516 6964 2524
rect 6956 2496 6964 2504
rect 6972 2476 6980 2484
rect 6956 2356 6964 2364
rect 6940 2316 6948 2324
rect 6940 2296 6948 2304
rect 6892 2276 6900 2284
rect 6924 2256 6932 2264
rect 6924 2196 6932 2204
rect 6940 2176 6948 2184
rect 6892 2156 6900 2164
rect 6908 2136 6916 2144
rect 6876 2116 6884 2124
rect 6860 1916 6868 1924
rect 6812 1876 6820 1884
rect 6844 1876 6852 1884
rect 6860 1756 6868 1764
rect 6812 1736 6820 1744
rect 6828 1696 6836 1704
rect 6844 1536 6852 1544
rect 6780 1476 6788 1484
rect 6748 1436 6756 1444
rect 6780 1436 6788 1444
rect 6764 1396 6772 1404
rect 6732 1376 6740 1384
rect 6764 1356 6772 1364
rect 6796 1416 6804 1424
rect 6972 2336 6980 2344
rect 6972 2236 6980 2244
rect 6988 2156 6996 2164
rect 6940 1916 6948 1924
rect 6956 1916 6964 1924
rect 6892 1896 6900 1904
rect 6892 1876 6900 1884
rect 6908 1856 6916 1864
rect 6956 1896 6964 1904
rect 6956 1856 6964 1864
rect 6924 1816 6932 1824
rect 6924 1756 6932 1764
rect 6892 1716 6900 1724
rect 6924 1676 6932 1684
rect 6876 1536 6884 1544
rect 6940 1536 6948 1544
rect 6988 1816 6996 1824
rect 6972 1736 6980 1744
rect 7180 3756 7188 3764
rect 7196 3736 7204 3744
rect 7100 3676 7108 3684
rect 7132 3716 7140 3724
rect 7164 3656 7172 3664
rect 7116 3636 7124 3644
rect 7116 3616 7124 3624
rect 7308 4296 7316 4304
rect 7276 4016 7284 4024
rect 7228 3896 7236 3904
rect 7276 3896 7284 3904
rect 7260 3876 7268 3884
rect 7292 3856 7300 3864
rect 7260 3836 7268 3844
rect 7228 3756 7236 3764
rect 7180 3576 7188 3584
rect 7180 3536 7188 3544
rect 7132 3516 7140 3524
rect 7212 3556 7220 3564
rect 7164 3496 7172 3504
rect 7132 3476 7140 3484
rect 7116 3416 7124 3424
rect 7132 3376 7140 3384
rect 7244 3476 7252 3484
rect 7340 3756 7348 3764
rect 7276 3716 7284 3724
rect 7324 3716 7332 3724
rect 7292 3496 7300 3504
rect 7212 3376 7220 3384
rect 7148 3356 7156 3364
rect 7164 3356 7172 3364
rect 7212 3356 7220 3364
rect 7164 3336 7172 3344
rect 7180 3316 7188 3324
rect 7116 3296 7124 3304
rect 7100 3256 7108 3264
rect 7164 3256 7172 3264
rect 7132 3216 7140 3224
rect 7116 3136 7124 3144
rect 7084 3056 7092 3064
rect 7052 3036 7060 3044
rect 7068 2936 7076 2944
rect 7052 2916 7060 2924
rect 7068 2716 7076 2724
rect 7084 2716 7092 2724
rect 7052 2616 7060 2624
rect 7036 2596 7044 2604
rect 7116 2896 7124 2904
rect 7116 2656 7124 2664
rect 7100 2576 7108 2584
rect 7148 3176 7156 3184
rect 7196 3276 7204 3284
rect 7164 2916 7172 2924
rect 7180 2836 7188 2844
rect 7164 2676 7172 2684
rect 7196 2676 7204 2684
rect 7132 2616 7140 2624
rect 7148 2576 7156 2584
rect 7180 2576 7188 2584
rect 7100 2496 7108 2504
rect 7116 2276 7124 2284
rect 7100 2216 7108 2224
rect 7132 2216 7140 2224
rect 7084 2136 7092 2144
rect 7116 2136 7124 2144
rect 7036 2116 7044 2124
rect 7052 2116 7060 2124
rect 7084 2116 7092 2124
rect 7052 2076 7060 2084
rect 7068 1896 7076 1904
rect 7052 1856 7060 1864
rect 7036 1796 7044 1804
rect 7036 1736 7044 1744
rect 6972 1716 6980 1724
rect 7036 1716 7044 1724
rect 7020 1576 7028 1584
rect 6988 1536 6996 1544
rect 6956 1496 6964 1504
rect 6876 1476 6884 1484
rect 6860 1416 6868 1424
rect 6812 1336 6820 1344
rect 6844 1336 6852 1344
rect 6716 1296 6724 1304
rect 6748 1276 6756 1284
rect 6732 1076 6740 1084
rect 6700 1056 6708 1064
rect 6764 976 6772 984
rect 6668 956 6676 964
rect 6748 956 6756 964
rect 6844 1276 6852 1284
rect 6860 1236 6868 1244
rect 6796 1176 6804 1184
rect 6684 936 6692 944
rect 6780 936 6788 944
rect 6828 1076 6836 1084
rect 6924 1476 6932 1484
rect 6908 1416 6916 1424
rect 6892 1396 6900 1404
rect 6988 1496 6996 1504
rect 6988 1456 6996 1464
rect 6892 1316 6900 1324
rect 6892 1296 6900 1304
rect 6924 1276 6932 1284
rect 6908 1216 6916 1224
rect 6972 1136 6980 1144
rect 6972 1116 6980 1124
rect 6956 1096 6964 1104
rect 6876 956 6884 964
rect 6908 936 6916 944
rect 6700 756 6708 764
rect 6684 736 6692 744
rect 6812 916 6820 924
rect 6892 916 6900 924
rect 6796 856 6804 864
rect 6796 796 6804 804
rect 6892 896 6900 904
rect 6828 836 6836 844
rect 6844 776 6852 784
rect 6812 736 6820 744
rect 6860 736 6868 744
rect 6716 716 6724 724
rect 6732 696 6740 704
rect 6684 676 6692 684
rect 6780 676 6788 684
rect 6796 676 6804 684
rect 6748 656 6756 664
rect 6780 556 6788 564
rect 6828 696 6836 704
rect 6844 696 6852 704
rect 6812 656 6820 664
rect 6828 656 6836 664
rect 6876 596 6884 604
rect 6812 556 6820 564
rect 6748 536 6756 544
rect 6764 536 6772 544
rect 6844 536 6852 544
rect 6684 516 6692 524
rect 6860 516 6868 524
rect 6732 336 6740 344
rect 6828 336 6836 344
rect 6732 316 6740 324
rect 6844 316 6852 324
rect 6700 276 6708 284
rect 6716 236 6724 244
rect 6924 836 6932 844
rect 6940 816 6948 824
rect 7004 1396 7012 1404
rect 7052 1676 7060 1684
rect 7116 2096 7124 2104
rect 7180 2396 7188 2404
rect 7164 2216 7172 2224
rect 7148 2116 7156 2124
rect 7100 1916 7108 1924
rect 7116 1876 7124 1884
rect 7100 1856 7108 1864
rect 7084 1736 7092 1744
rect 7084 1716 7092 1724
rect 7068 1576 7076 1584
rect 7052 1556 7060 1564
rect 7084 1536 7092 1544
rect 7036 1496 7044 1504
rect 7052 1496 7060 1504
rect 7084 1456 7092 1464
rect 7068 1416 7076 1424
rect 7164 2076 7172 2084
rect 7164 2036 7172 2044
rect 7372 3716 7380 3724
rect 7372 3516 7380 3524
rect 7292 3336 7300 3344
rect 7308 3336 7316 3344
rect 7276 3316 7284 3324
rect 7276 3276 7284 3284
rect 7244 3216 7252 3224
rect 7260 3156 7268 3164
rect 7308 3296 7316 3304
rect 7308 3076 7316 3084
rect 7356 3236 7364 3244
rect 7340 3156 7348 3164
rect 7340 3076 7348 3084
rect 7244 2936 7252 2944
rect 7244 2676 7252 2684
rect 7260 2436 7268 2444
rect 7196 2176 7204 2184
rect 7180 2016 7188 2024
rect 7180 1996 7188 2004
rect 7180 1856 7188 1864
rect 7228 1996 7236 2004
rect 7244 1876 7252 1884
rect 7148 1836 7156 1844
rect 7196 1836 7204 1844
rect 7180 1816 7188 1824
rect 7132 1776 7140 1784
rect 7164 1756 7172 1764
rect 7148 1736 7156 1744
rect 7132 1716 7140 1724
rect 7132 1696 7140 1704
rect 7164 1676 7172 1684
rect 7180 1656 7188 1664
rect 7148 1616 7156 1624
rect 7180 1616 7188 1624
rect 7212 1596 7220 1604
rect 7196 1576 7204 1584
rect 7196 1536 7204 1544
rect 7100 1396 7108 1404
rect 7116 1356 7124 1364
rect 7036 1336 7044 1344
rect 7132 1336 7140 1344
rect 7036 1296 7044 1304
rect 7020 1156 7028 1164
rect 7084 1156 7092 1164
rect 7020 1056 7028 1064
rect 6988 936 6996 944
rect 6988 916 6996 924
rect 7052 916 7060 924
rect 6972 896 6980 904
rect 7004 896 7012 904
rect 6988 876 6996 884
rect 6956 756 6964 764
rect 7004 756 7012 764
rect 6908 736 6916 744
rect 6956 736 6964 744
rect 6908 716 6916 724
rect 6956 696 6964 704
rect 6924 676 6932 684
rect 6956 676 6964 684
rect 6908 576 6916 584
rect 6924 556 6932 564
rect 6892 536 6900 544
rect 6892 496 6900 504
rect 6972 596 6980 604
rect 7068 696 7076 704
rect 7020 676 7028 684
rect 7052 576 7060 584
rect 7052 516 7060 524
rect 7036 496 7044 504
rect 7004 436 7012 444
rect 6972 316 6980 324
rect 7004 296 7012 304
rect 7036 276 7044 284
rect 6876 256 6884 264
rect 6860 216 6868 224
rect 6620 196 6628 204
rect 6652 196 6660 204
rect 6812 196 6820 204
rect 6684 176 6692 184
rect 6892 156 6900 164
rect 6940 156 6948 164
rect 7052 176 7060 184
rect 7116 1136 7124 1144
rect 7100 1076 7108 1084
rect 7116 656 7124 664
rect 7100 616 7108 624
rect 7116 576 7124 584
rect 7116 536 7124 544
rect 7164 1476 7172 1484
rect 7180 1436 7188 1444
rect 7148 1316 7156 1324
rect 7324 2816 7332 2824
rect 7340 2716 7348 2724
rect 7356 2696 7364 2704
rect 7404 3316 7412 3324
rect 7388 3016 7396 3024
rect 7404 2756 7412 2764
rect 7292 2516 7300 2524
rect 7308 2302 7316 2304
rect 7308 2296 7316 2302
rect 7372 2576 7380 2584
rect 7340 2176 7348 2184
rect 7292 2096 7300 2104
rect 7276 1856 7284 1864
rect 7276 1836 7284 1844
rect 7276 1756 7284 1764
rect 7276 1696 7284 1704
rect 7276 1556 7284 1564
rect 7228 1536 7236 1544
rect 7228 1496 7236 1504
rect 7244 1476 7252 1484
rect 7164 976 7172 984
rect 7148 696 7156 704
rect 7148 596 7156 604
rect 7228 1316 7236 1324
rect 7244 1116 7252 1124
rect 7228 1076 7236 1084
rect 7228 976 7236 984
rect 7260 1076 7268 1084
rect 7260 1056 7268 1064
rect 7244 956 7252 964
rect 7212 916 7220 924
rect 7244 916 7252 924
rect 7260 916 7268 924
rect 7244 896 7252 904
rect 7228 876 7236 884
rect 7228 736 7236 744
rect 7212 696 7220 704
rect 7212 676 7220 684
rect 7196 656 7204 664
rect 7148 556 7156 564
rect 7180 576 7188 584
rect 7340 2016 7348 2024
rect 7308 1902 7316 1904
rect 7308 1896 7316 1902
rect 7356 1836 7364 1844
rect 7324 1776 7332 1784
rect 7340 1776 7348 1784
rect 7292 1476 7300 1484
rect 7372 1816 7380 1824
rect 7356 1536 7364 1544
rect 7340 1516 7348 1524
rect 7340 1396 7348 1404
rect 7308 1336 7316 1344
rect 7292 1116 7300 1124
rect 7292 1016 7300 1024
rect 7372 1096 7380 1104
rect 7324 1076 7332 1084
rect 7356 1056 7364 1064
rect 7308 996 7316 1004
rect 7356 1036 7364 1044
rect 7276 876 7284 884
rect 7260 816 7268 824
rect 7340 976 7348 984
rect 7340 936 7348 944
rect 7308 916 7316 924
rect 7292 796 7300 804
rect 7308 696 7316 704
rect 7244 556 7252 564
rect 7244 516 7252 524
rect 7276 656 7284 664
rect 7372 956 7380 964
rect 7356 816 7364 824
rect 7356 796 7364 804
rect 7340 656 7348 664
rect 7324 636 7332 644
rect 7292 616 7300 624
rect 7260 356 7268 364
rect 7260 296 7268 304
rect 7164 276 7172 284
rect 7196 276 7204 284
rect 7404 1796 7412 1804
rect 7388 196 7396 204
rect 7084 156 7092 164
rect 7036 136 7044 144
rect 7196 136 7204 144
rect 7340 136 7348 144
rect 6844 116 6852 124
rect 7212 116 7220 124
rect 6044 96 6052 104
rect 6156 96 6164 104
rect 6652 96 6660 104
rect 7068 96 7076 104
rect 5196 16 5204 24
<< metal3 >>
rect 2564 5417 2588 5423
rect 3476 5417 3500 5423
rect 3620 5417 3644 5423
rect 2914 5414 2974 5416
rect 2914 5406 2915 5414
rect 2924 5406 2925 5414
rect 2963 5406 2964 5414
rect 2973 5406 2974 5414
rect 2914 5404 2974 5406
rect 5922 5414 5982 5416
rect 5922 5406 5923 5414
rect 5932 5406 5933 5414
rect 5971 5406 5972 5414
rect 5981 5406 5982 5414
rect 5922 5404 5982 5406
rect 1044 5397 1100 5403
rect 3444 5397 3468 5403
rect 4324 5397 5644 5403
rect 6932 5397 7052 5403
rect 468 5377 508 5383
rect 797 5377 1324 5383
rect 797 5364 803 5377
rect 1332 5377 1484 5383
rect 1924 5377 2028 5383
rect 2292 5377 2332 5383
rect 3364 5377 3452 5383
rect 3732 5377 3916 5383
rect 3924 5377 4396 5383
rect 4404 5377 4556 5383
rect 5444 5377 5628 5383
rect 5764 5377 5852 5383
rect 5860 5377 6492 5383
rect 6500 5377 6604 5383
rect 6804 5377 6988 5383
rect 324 5357 396 5363
rect 404 5357 620 5363
rect 628 5357 796 5363
rect 852 5357 956 5363
rect 1092 5357 1212 5363
rect 1220 5357 1276 5363
rect 1284 5357 1564 5363
rect 1572 5357 1644 5363
rect 1652 5357 1836 5363
rect 1908 5357 1964 5363
rect 2004 5357 2076 5363
rect 2084 5357 2108 5363
rect 2212 5357 2380 5363
rect 2388 5357 2684 5363
rect 3076 5357 3404 5363
rect 4212 5357 4316 5363
rect 5300 5357 5324 5363
rect 5348 5357 5420 5363
rect 5572 5357 5676 5363
rect 5812 5357 5900 5363
rect 5908 5357 5996 5363
rect 6004 5357 6188 5363
rect 6324 5357 6412 5363
rect 6420 5357 7196 5363
rect 292 5337 364 5343
rect 388 5337 428 5343
rect 436 5337 492 5343
rect 500 5337 540 5343
rect 548 5337 572 5343
rect 580 5337 748 5343
rect 772 5337 796 5343
rect 893 5337 1068 5343
rect 52 5317 156 5323
rect 212 5317 652 5323
rect 708 5317 764 5323
rect 893 5323 899 5337
rect 1604 5337 1612 5343
rect 1636 5337 1692 5343
rect 1821 5337 2524 5343
rect 772 5317 899 5323
rect 916 5317 1004 5323
rect 1012 5317 1052 5323
rect 1821 5323 1827 5337
rect 2532 5337 2588 5343
rect 2756 5337 3100 5343
rect 3108 5337 3212 5343
rect 3348 5337 3420 5343
rect 3428 5337 3468 5343
rect 3476 5337 3548 5343
rect 3860 5337 3948 5343
rect 4660 5337 4796 5343
rect 5268 5337 5596 5343
rect 5604 5337 6060 5343
rect 6132 5337 6220 5343
rect 6372 5337 6460 5343
rect 6468 5337 6796 5343
rect 7021 5337 7068 5343
rect 7021 5324 7027 5337
rect 1188 5317 1827 5323
rect 1860 5317 1916 5323
rect 1940 5317 2044 5323
rect 2052 5317 2204 5323
rect 2276 5317 2316 5323
rect 2372 5317 2428 5323
rect 2724 5317 3500 5323
rect 3572 5317 4035 5323
rect -35 5297 12 5303
rect 116 5297 1180 5303
rect 1508 5297 1596 5303
rect 1604 5297 1660 5303
rect 1684 5297 1788 5303
rect 1812 5297 1932 5303
rect 1988 5297 2092 5303
rect 2100 5297 2220 5303
rect 2532 5297 2556 5303
rect 2692 5297 3212 5303
rect 3220 5297 3324 5303
rect 3380 5297 3484 5303
rect 3572 5297 3596 5303
rect 3956 5297 3996 5303
rect 4004 5297 4012 5303
rect 4029 5303 4035 5317
rect 4116 5317 4252 5323
rect 4356 5317 4508 5323
rect 4516 5317 4588 5323
rect 4596 5317 4700 5323
rect 4836 5317 4972 5323
rect 5060 5317 5196 5323
rect 5316 5317 5324 5323
rect 5668 5317 5708 5323
rect 6228 5317 6268 5323
rect 6276 5317 7020 5323
rect 7172 5317 7308 5323
rect 4029 5297 4924 5303
rect 4964 5297 5308 5303
rect 5364 5297 5372 5303
rect 5428 5297 5772 5303
rect 5828 5297 6364 5303
rect 6532 5297 6572 5303
rect 6580 5297 7100 5303
rect 7108 5297 7164 5303
rect 7204 5297 7276 5303
rect 660 5277 2172 5283
rect 2180 5277 2940 5283
rect 3460 5277 5372 5283
rect 5636 5277 5852 5283
rect 6484 5277 6540 5283
rect 6580 5277 6716 5283
rect 260 5257 668 5263
rect 756 5257 844 5263
rect 852 5257 892 5263
rect 980 5257 1132 5263
rect 1140 5257 1356 5263
rect 1364 5257 1612 5263
rect 1700 5257 2092 5263
rect 2100 5257 2156 5263
rect 4244 5257 4300 5263
rect 4628 5257 4668 5263
rect 4676 5257 5804 5263
rect 5908 5257 6428 5263
rect 820 5237 1020 5243
rect 1028 5237 1372 5243
rect 1380 5237 1404 5243
rect 1716 5237 1756 5243
rect 1764 5237 2012 5243
rect 3428 5237 3468 5243
rect 4212 5237 4988 5243
rect 4996 5237 5452 5243
rect 5460 5237 6572 5243
rect 6580 5237 7004 5243
rect 7012 5237 7084 5243
rect 324 5217 1164 5223
rect 2788 5217 2988 5223
rect 4644 5217 5004 5223
rect 5012 5217 5052 5223
rect 5060 5217 5660 5223
rect 5732 5217 6284 5223
rect 6292 5217 6588 5223
rect 6596 5217 7276 5223
rect 1410 5214 1470 5216
rect 1410 5206 1411 5214
rect 1420 5206 1421 5214
rect 1459 5206 1460 5214
rect 1469 5206 1470 5214
rect 1410 5204 1470 5206
rect 4418 5214 4478 5216
rect 4418 5206 4419 5214
rect 4428 5206 4429 5214
rect 4467 5206 4468 5214
rect 4477 5206 4478 5214
rect 4418 5204 4478 5206
rect 1828 5197 2108 5203
rect 2276 5197 2780 5203
rect 4916 5197 5020 5203
rect 5348 5197 6124 5203
rect 868 5177 1116 5183
rect 1332 5177 1804 5183
rect 1828 5177 1900 5183
rect 1908 5177 1916 5183
rect 2020 5177 2044 5183
rect 2052 5177 2268 5183
rect 2372 5177 2668 5183
rect 4548 5177 4796 5183
rect 5092 5177 5484 5183
rect 5588 5177 6332 5183
rect 1108 5157 1148 5163
rect 1172 5157 1868 5163
rect 1876 5157 2796 5163
rect 2804 5157 3132 5163
rect 4580 5157 5116 5163
rect 5124 5157 5196 5163
rect 5204 5157 5404 5163
rect 5412 5157 5500 5163
rect 5508 5157 5996 5163
rect 6164 5157 6332 5163
rect 980 5137 1164 5143
rect 1236 5137 1436 5143
rect 1492 5137 1596 5143
rect 1844 5137 1932 5143
rect 2212 5137 2476 5143
rect 2484 5137 2924 5143
rect 2932 5137 3260 5143
rect 3268 5137 3436 5143
rect 4692 5137 4716 5143
rect 5316 5137 5356 5143
rect 5380 5137 5740 5143
rect 5812 5137 5884 5143
rect 6020 5137 6156 5143
rect 6164 5137 6988 5143
rect 6996 5137 7180 5143
rect 532 5117 556 5123
rect 612 5117 636 5123
rect 692 5117 2243 5123
rect 2237 5104 2243 5117
rect 2292 5117 2348 5123
rect 2436 5117 2460 5123
rect 2845 5117 3052 5123
rect 2845 5104 2851 5117
rect 3220 5117 3308 5123
rect 3364 5117 3484 5123
rect 3492 5117 3596 5123
rect 4020 5117 4236 5123
rect 4388 5117 4620 5123
rect 4660 5117 4748 5123
rect 4900 5117 5148 5123
rect 5172 5117 5228 5123
rect 5252 5117 5324 5123
rect 5332 5117 5436 5123
rect 5716 5117 5724 5123
rect 5844 5117 5868 5123
rect 6228 5117 6300 5123
rect 6468 5117 6636 5123
rect 7124 5117 7228 5123
rect 20 5097 60 5103
rect 116 5097 156 5103
rect 164 5097 188 5103
rect 212 5097 236 5103
rect 308 5097 332 5103
rect 340 5097 380 5103
rect 420 5097 556 5103
rect 596 5097 636 5103
rect 644 5097 748 5103
rect 756 5097 796 5103
rect 804 5097 828 5103
rect 964 5097 1036 5103
rect 1060 5097 1100 5103
rect 1108 5097 1148 5103
rect 1172 5097 1196 5103
rect 1220 5097 1260 5103
rect 1316 5097 1324 5103
rect 1524 5097 1548 5103
rect 1556 5097 1660 5103
rect 1796 5097 1836 5103
rect 2244 5097 2844 5103
rect 2900 5097 3244 5103
rect 3380 5097 3484 5103
rect 3540 5097 3564 5103
rect 3748 5097 3964 5103
rect 4116 5097 4268 5103
rect 4340 5097 4707 5103
rect 189 5083 195 5096
rect 189 5077 236 5083
rect 404 5077 444 5083
rect 548 5077 716 5083
rect 724 5077 812 5083
rect 1012 5077 1036 5083
rect 1140 5077 1212 5083
rect 1220 5077 1692 5083
rect 1700 5077 1708 5083
rect 1716 5077 1724 5083
rect 1732 5077 1804 5083
rect 1860 5077 1939 5083
rect 84 5057 124 5063
rect 132 5057 220 5063
rect 228 5057 252 5063
rect 260 5057 300 5063
rect 436 5057 492 5063
rect 676 5057 732 5063
rect 740 5057 828 5063
rect 836 5057 892 5063
rect 900 5057 1020 5063
rect 1300 5057 1340 5063
rect 1348 5057 1676 5063
rect 1684 5057 1692 5063
rect 1700 5057 1900 5063
rect 1933 5063 1939 5077
rect 2116 5077 2156 5083
rect 2308 5077 2380 5083
rect 2452 5077 2604 5083
rect 2820 5077 2876 5083
rect 3460 5077 3532 5083
rect 3988 5077 4284 5083
rect 4372 5077 4460 5083
rect 4612 5077 4652 5083
rect 4701 5083 4707 5097
rect 4772 5097 5420 5103
rect 5428 5097 5548 5103
rect 5892 5097 5916 5103
rect 5924 5097 6172 5103
rect 6196 5097 6268 5103
rect 6564 5097 6716 5103
rect 6772 5097 6828 5103
rect 6868 5097 7308 5103
rect 4701 5077 4860 5083
rect 4868 5077 4908 5083
rect 5012 5077 5084 5083
rect 5172 5077 5212 5083
rect 5220 5077 5468 5083
rect 5476 5077 5484 5083
rect 5556 5077 5628 5083
rect 5645 5077 5820 5083
rect 1933 5057 2108 5063
rect 2116 5057 2540 5063
rect 2548 5057 3180 5063
rect 4260 5057 4300 5063
rect 4308 5057 4556 5063
rect 4564 5057 5260 5063
rect 5316 5057 5340 5063
rect 5645 5063 5651 5077
rect 6276 5077 6524 5083
rect 6532 5077 6572 5083
rect 6644 5077 6908 5083
rect 6964 5077 7148 5083
rect 7156 5077 7196 5083
rect 7220 5077 7260 5083
rect 7300 5077 7372 5083
rect 5412 5057 5651 5063
rect 5684 5057 5724 5063
rect 5748 5057 6028 5063
rect 6116 5057 6220 5063
rect 6260 5057 6412 5063
rect 84 5037 348 5043
rect 868 5037 1644 5043
rect 1652 5037 2268 5043
rect 2276 5037 3516 5043
rect 3524 5037 3612 5043
rect 4052 5037 4204 5043
rect 4228 5037 4332 5043
rect 4436 5037 4588 5043
rect 4596 5037 4620 5043
rect 4628 5037 4684 5043
rect 4708 5037 4876 5043
rect 5076 5037 5132 5043
rect 5140 5037 5196 5043
rect 5213 5037 5372 5043
rect 500 5017 972 5023
rect 1012 5017 1068 5023
rect 1780 5017 1868 5023
rect 1876 5017 1996 5023
rect 2052 5017 2563 5023
rect 532 4997 604 5003
rect 1252 4997 1356 5003
rect 1764 4997 2172 5003
rect 2180 4997 2220 5003
rect 2340 4997 2540 5003
rect 2557 5003 2563 5017
rect 2580 5017 2588 5023
rect 2788 5017 2892 5023
rect 3236 5017 3356 5023
rect 3556 5017 4716 5023
rect 4740 5017 4844 5023
rect 5213 5023 5219 5037
rect 5444 5037 5740 5043
rect 5812 5037 5852 5043
rect 5860 5037 5932 5043
rect 6180 5037 6268 5043
rect 6500 5037 6604 5043
rect 7108 5037 7116 5043
rect 7316 5037 7340 5043
rect 5060 5017 5219 5023
rect 5332 5017 5708 5023
rect 5796 5017 5900 5023
rect 6388 5017 6460 5023
rect 2914 5014 2974 5016
rect 2914 5006 2915 5014
rect 2924 5006 2925 5014
rect 2963 5006 2964 5014
rect 2973 5006 2974 5014
rect 2914 5004 2974 5006
rect 5922 5014 5982 5016
rect 5922 5006 5923 5014
rect 5932 5006 5933 5014
rect 5971 5006 5972 5014
rect 5981 5006 5982 5014
rect 5922 5004 5982 5006
rect 2557 4997 2636 5003
rect 3044 4997 3100 5003
rect 3284 4997 3388 5003
rect 4020 4997 4572 5003
rect 4612 4997 4620 5003
rect 4756 4997 4796 5003
rect 4820 4997 4860 5003
rect 4964 4997 5116 5003
rect 5124 4997 5692 5003
rect 5700 4997 5852 5003
rect 6084 4997 6211 5003
rect 68 4977 108 4983
rect 212 4977 252 4983
rect 404 4977 684 4983
rect 1300 4977 1308 4983
rect 1316 4977 1516 4983
rect 1828 4977 2028 4983
rect 2084 4977 2412 4983
rect 2500 4977 2620 4983
rect 2733 4977 3580 4983
rect 2733 4964 2739 4977
rect 4260 4977 4444 4983
rect 4452 4977 4988 4983
rect 4996 4977 5180 4983
rect 5428 4977 5555 4983
rect 5549 4964 5555 4977
rect 5652 4977 5715 4983
rect 212 4957 332 4963
rect 548 4957 588 4963
rect 612 4957 684 4963
rect 724 4957 908 4963
rect 996 4957 1148 4963
rect 1236 4957 1260 4963
rect 1284 4957 1420 4963
rect 1444 4957 1500 4963
rect 1508 4957 1532 4963
rect 1540 4957 1580 4963
rect 1620 4957 1795 4963
rect 148 4937 252 4943
rect 500 4937 508 4943
rect 516 4937 588 4943
rect 628 4937 668 4943
rect 676 4937 940 4943
rect 948 4937 988 4943
rect 996 4937 1068 4943
rect 1172 4937 1196 4943
rect 1284 4937 1372 4943
rect 1524 4937 1580 4943
rect 1789 4943 1795 4957
rect 1812 4957 1852 4963
rect 1972 4957 2076 4963
rect 2260 4957 2300 4963
rect 2372 4957 2460 4963
rect 2468 4957 2732 4963
rect 2836 4957 3084 4963
rect 3092 4957 3292 4963
rect 3684 4957 3788 4963
rect 4148 4957 4556 4963
rect 4580 4957 4764 4963
rect 5028 4957 5068 4963
rect 5108 4957 5164 4963
rect 5364 4957 5516 4963
rect 5556 4957 5644 4963
rect 5652 4957 5692 4963
rect 5709 4963 5715 4977
rect 5892 4977 6188 4983
rect 6205 4983 6211 4997
rect 6292 4997 6348 5003
rect 6356 4997 6556 5003
rect 6564 4997 6796 5003
rect 6205 4977 6396 4983
rect 6436 4977 6524 4983
rect 6532 4977 6940 4983
rect 6948 4977 7180 4983
rect 5709 4957 6012 4963
rect 6020 4957 6140 4963
rect 6212 4957 6460 4963
rect 6596 4957 6652 4963
rect 6916 4957 6988 4963
rect 6996 4957 7100 4963
rect 7108 4957 7212 4963
rect 1789 4937 1836 4943
rect 1876 4937 1996 4943
rect 2164 4937 2252 4943
rect 2484 4937 2508 4943
rect 2532 4937 2588 4943
rect 2900 4937 3052 4943
rect 3412 4937 3468 4943
rect 3540 4937 3676 4943
rect 3924 4937 3964 4943
rect 4052 4937 4060 4943
rect 4244 4937 4332 4943
rect 4356 4937 4396 4943
rect 4916 4937 5068 4943
rect 5101 4937 5132 4943
rect 180 4917 220 4923
rect 372 4917 412 4923
rect 580 4917 732 4923
rect 948 4917 972 4923
rect 980 4917 1004 4923
rect 1044 4917 1116 4923
rect 1252 4917 1260 4923
rect 1332 4917 1596 4923
rect 1764 4917 1772 4923
rect 1780 4917 1964 4923
rect 1988 4917 2060 4923
rect 2100 4917 2124 4923
rect 2164 4917 2236 4923
rect 2420 4917 2476 4923
rect 2724 4917 2803 4923
rect -35 4897 316 4903
rect 772 4897 924 4903
rect 932 4897 1324 4903
rect 1332 4897 2780 4903
rect 2797 4903 2803 4917
rect 3204 4917 3276 4923
rect 3284 4917 3324 4923
rect 3332 4917 3404 4923
rect 3540 4917 3580 4923
rect 3668 4917 3820 4923
rect 4628 4917 4876 4923
rect 5101 4923 5107 4937
rect 5140 4937 5388 4943
rect 5428 4937 5612 4943
rect 5732 4937 5756 4943
rect 5812 4937 6172 4943
rect 6180 4937 6220 4943
rect 6340 4937 6364 4943
rect 6372 4937 6444 4943
rect 6452 4937 6668 4943
rect 6692 4937 6780 4943
rect 6788 4937 6956 4943
rect 6964 4937 7052 4943
rect 4884 4917 5107 4923
rect 5124 4917 5260 4923
rect 5316 4917 5468 4923
rect 5716 4917 5724 4923
rect 5748 4917 5772 4923
rect 5860 4917 5964 4923
rect 6036 4917 6300 4923
rect 6388 4917 6476 4923
rect 6740 4917 6828 4923
rect 6980 4917 7292 4923
rect 2797 4897 3244 4903
rect 3604 4897 3628 4903
rect 3636 4897 3900 4903
rect 4548 4897 4604 4903
rect 4660 4897 5100 4903
rect 5220 4897 5596 4903
rect 5796 4897 5836 4903
rect 6036 4897 6860 4903
rect 7124 4897 7132 4903
rect 484 4877 636 4883
rect 1268 4877 1324 4883
rect 1348 4877 1372 4883
rect 1380 4877 2428 4883
rect 3060 4877 3132 4883
rect 3172 4877 3260 4883
rect 3268 4877 3484 4883
rect 3700 4877 5868 4883
rect 6164 4877 6268 4883
rect 1364 4857 1404 4863
rect 1428 4857 1980 4863
rect 2068 4857 2316 4863
rect 2564 4857 2604 4863
rect 2628 4857 2924 4863
rect 2932 4857 3340 4863
rect 3348 4857 3388 4863
rect 3485 4863 3491 4876
rect 3485 4857 3948 4863
rect 4196 4857 4492 4863
rect 4596 4857 4684 4863
rect 4740 4857 4764 4863
rect 5012 4857 5036 4863
rect 5092 4857 5116 4863
rect 5124 4857 5564 4863
rect 5588 4857 5692 4863
rect 5764 4857 6092 4863
rect 6100 4857 6300 4863
rect 6308 4857 6412 4863
rect 980 4837 1532 4843
rect 1668 4837 1836 4843
rect 1876 4837 2332 4843
rect 2420 4837 2460 4843
rect 2516 4837 2572 4843
rect 2580 4837 2988 4843
rect 3092 4837 3164 4843
rect 3220 4837 3292 4843
rect 3460 4837 3468 4843
rect 3860 4837 3932 4843
rect 3940 4837 3996 4843
rect 4004 4837 4076 4843
rect 4324 4837 5331 4843
rect 1620 4817 1932 4823
rect 2084 4817 2604 4823
rect 3348 4817 3868 4823
rect 4532 4817 4652 4823
rect 4676 4817 5308 4823
rect 5325 4823 5331 4837
rect 5364 4837 5756 4843
rect 5796 4837 5804 4843
rect 5812 4837 6188 4843
rect 6212 4837 6284 4843
rect 6292 4837 6540 4843
rect 6548 4837 6764 4843
rect 5325 4817 5596 4823
rect 5620 4817 6044 4823
rect 6068 4817 6108 4823
rect 1410 4814 1470 4816
rect 1410 4806 1411 4814
rect 1420 4806 1421 4814
rect 1459 4806 1460 4814
rect 1469 4806 1470 4814
rect 1410 4804 1470 4806
rect 4418 4814 4478 4816
rect 4418 4806 4419 4814
rect 4428 4806 4429 4814
rect 4467 4806 4468 4814
rect 4477 4806 4478 4814
rect 4418 4804 4478 4806
rect 436 4797 1395 4803
rect 1389 4783 1395 4797
rect 2212 4797 2428 4803
rect 2436 4797 2492 4803
rect 2516 4797 2700 4803
rect 3044 4797 3452 4803
rect 3572 4797 3628 4803
rect 3636 4797 3804 4803
rect 4532 4797 5916 4803
rect 6148 4797 6796 4803
rect 1108 4777 1315 4783
rect 1389 4777 1468 4783
rect 244 4757 508 4763
rect 516 4757 556 4763
rect 564 4757 588 4763
rect 989 4757 1052 4763
rect 989 4744 995 4757
rect 1060 4757 1100 4763
rect 1309 4763 1315 4777
rect 2308 4777 2604 4783
rect 2868 4777 3420 4783
rect 3444 4777 3500 4783
rect 3549 4777 3708 4783
rect 1309 4757 1676 4763
rect 1684 4757 2572 4763
rect 3549 4763 3555 4777
rect 4516 4777 4620 4783
rect 4628 4777 5164 4783
rect 5492 4777 5580 4783
rect 5604 4777 6268 4783
rect 6836 4777 6860 4783
rect 6868 4777 6972 4783
rect 2708 4757 3555 4763
rect 3572 4757 4524 4763
rect 4628 4757 4732 4763
rect 4740 4757 4780 4763
rect 4820 4757 5132 4763
rect 5172 4757 5420 4763
rect 5492 4757 5564 4763
rect 5668 4757 5788 4763
rect 5812 4757 5868 4763
rect 5908 4757 6108 4763
rect 6388 4757 6700 4763
rect 20 4737 44 4743
rect 52 4737 124 4743
rect 132 4737 140 4743
rect 148 4737 204 4743
rect 212 4737 364 4743
rect 740 4737 988 4743
rect 1060 4737 1116 4743
rect 1332 4737 1356 4743
rect 1588 4737 2012 4743
rect 2068 4737 2140 4743
rect 2212 4737 2540 4743
rect 2676 4737 2844 4743
rect 3316 4737 4108 4743
rect 4372 4737 4524 4743
rect 4644 4737 4700 4743
rect 4820 4737 5148 4743
rect 5156 4737 5516 4743
rect 5524 4737 5740 4743
rect 5780 4737 6652 4743
rect 164 4717 460 4723
rect 804 4717 844 4723
rect 900 4717 1004 4723
rect 1092 4717 1308 4723
rect 1316 4717 1356 4723
rect 1972 4717 2108 4723
rect 2372 4717 2572 4723
rect 4116 4717 4236 4723
rect 4500 4717 4844 4723
rect 4884 4717 4956 4723
rect 5092 4717 5180 4723
rect 5204 4717 5212 4723
rect 5220 4717 5372 4723
rect 5556 4717 5820 4723
rect 5828 4717 5964 4723
rect 6068 4717 6332 4723
rect 6356 4717 6428 4723
rect 6484 4717 6588 4723
rect 292 4697 332 4703
rect 340 4697 428 4703
rect 580 4697 620 4703
rect 628 4697 844 4703
rect 884 4697 1260 4703
rect 1284 4697 1372 4703
rect 1620 4697 1644 4703
rect 1732 4697 1788 4703
rect 1844 4697 1996 4703
rect 2004 4697 2028 4703
rect 2100 4697 2220 4703
rect 2292 4697 2300 4703
rect 2324 4697 2396 4703
rect 2772 4697 2828 4703
rect 2884 4697 3068 4703
rect 3396 4697 3596 4703
rect 4004 4697 4124 4703
rect 4157 4697 4204 4703
rect 4157 4684 4163 4697
rect 4212 4697 4284 4703
rect 4292 4697 4300 4703
rect 4308 4697 4348 4703
rect 4516 4697 4652 4703
rect 4948 4697 4956 4703
rect 4964 4697 5452 4703
rect 5460 4697 5708 4703
rect 5716 4697 5868 4703
rect 5956 4697 5996 4703
rect 6068 4697 6076 4703
rect 6132 4697 6156 4703
rect 6260 4697 6364 4703
rect 6820 4697 6892 4703
rect 6948 4697 7132 4703
rect 7140 4697 7228 4703
rect 148 4677 156 4683
rect 164 4677 300 4683
rect 820 4677 956 4683
rect 964 4677 1100 4683
rect 1188 4677 1292 4683
rect 1524 4677 1756 4683
rect 1972 4677 2172 4683
rect 2420 4677 2540 4683
rect 2548 4677 2652 4683
rect 2740 4677 2780 4683
rect 2996 4677 3139 4683
rect 3133 4664 3139 4677
rect 3412 4677 3564 4683
rect 4084 4677 4156 4683
rect 4340 4677 4636 4683
rect 4644 4677 4684 4683
rect 4692 4677 4716 4683
rect 4724 4677 4940 4683
rect 5044 4677 5628 4683
rect 5636 4677 5804 4683
rect 6020 4677 6204 4683
rect 6228 4677 6476 4683
rect 6516 4677 6556 4683
rect 6564 4677 6620 4683
rect 6756 4677 6844 4683
rect 244 4657 284 4663
rect 468 4657 636 4663
rect 676 4657 812 4663
rect 916 4657 1116 4663
rect 1124 4657 1340 4663
rect 1348 4657 1388 4663
rect 1396 4657 1580 4663
rect 1780 4657 1804 4663
rect 1940 4657 1996 4663
rect 2164 4657 2380 4663
rect 2660 4657 2684 4663
rect 2724 4657 3004 4663
rect 3140 4657 3180 4663
rect 3396 4657 3692 4663
rect 3844 4657 4188 4663
rect 4244 4657 4316 4663
rect 4692 4657 4732 4663
rect 4756 4657 4780 4663
rect 4788 4657 5004 4663
rect 5012 4657 5068 4663
rect 5124 4657 5244 4663
rect 5252 4657 5324 4663
rect 5396 4657 5724 4663
rect 5748 4657 5788 4663
rect 6100 4657 6172 4663
rect 6308 4657 6396 4663
rect 6548 4657 6700 4663
rect 356 4637 508 4643
rect 948 4637 1004 4643
rect 1012 4637 1068 4643
rect 1604 4637 1660 4643
rect 1668 4637 1724 4643
rect 1732 4637 1852 4643
rect 1860 4637 2060 4643
rect 2068 4637 2076 4643
rect 2084 4637 2204 4643
rect 2372 4637 3212 4643
rect 3316 4637 3500 4643
rect 4180 4637 4524 4643
rect 4772 4637 4924 4643
rect 5117 4643 5123 4656
rect 4932 4637 5123 4643
rect 5300 4637 5628 4643
rect 5668 4637 6659 4643
rect 228 4617 396 4623
rect 500 4617 716 4623
rect 820 4617 1052 4623
rect 1316 4617 1948 4623
rect 1956 4617 2380 4623
rect 2628 4617 2732 4623
rect 2996 4617 3084 4623
rect 3213 4623 3219 4636
rect 3213 4617 3452 4623
rect 3460 4617 3580 4623
rect 3652 4617 3708 4623
rect 4020 4617 4972 4623
rect 4980 4617 5500 4623
rect 5508 4617 5548 4623
rect 5556 4617 5724 4623
rect 6004 4617 6140 4623
rect 6244 4617 6444 4623
rect 6452 4617 6476 4623
rect 6484 4617 6588 4623
rect 6653 4623 6659 4637
rect 6676 4637 7164 4643
rect 6653 4617 6748 4623
rect 6756 4617 6780 4623
rect 6932 4617 7084 4623
rect 2914 4614 2974 4616
rect 2914 4606 2915 4614
rect 2924 4606 2925 4614
rect 2963 4606 2964 4614
rect 2973 4606 2974 4614
rect 2914 4604 2974 4606
rect 5922 4614 5982 4616
rect 5922 4606 5923 4614
rect 5932 4606 5933 4614
rect 5971 4606 5972 4614
rect 5981 4606 5982 4614
rect 5922 4604 5982 4606
rect 644 4597 700 4603
rect 708 4597 764 4603
rect 1172 4597 1212 4603
rect 1572 4597 1756 4603
rect 1924 4597 1964 4603
rect 2468 4597 2556 4603
rect 2564 4597 2684 4603
rect 2692 4597 2876 4603
rect 2989 4597 3228 4603
rect 276 4577 316 4583
rect 340 4577 444 4583
rect 452 4577 476 4583
rect 724 4577 844 4583
rect 1028 4577 1084 4583
rect 1204 4577 1292 4583
rect 1988 4577 2156 4583
rect 2164 4577 2220 4583
rect 2244 4577 2316 4583
rect 2596 4577 2668 4583
rect 2733 4577 2764 4583
rect 84 4557 124 4563
rect 436 4557 492 4563
rect 500 4557 524 4563
rect 532 4557 588 4563
rect 836 4557 892 4563
rect 900 4557 924 4563
rect 932 4557 1132 4563
rect 1716 4557 1740 4563
rect 2084 4557 2140 4563
rect 2148 4557 2204 4563
rect 2324 4557 2380 4563
rect 2388 4557 2540 4563
rect 2733 4563 2739 4577
rect 2989 4583 2995 4597
rect 3412 4597 3436 4603
rect 3492 4597 3532 4603
rect 3588 4597 4691 4603
rect 2788 4577 2995 4583
rect 3172 4577 3548 4583
rect 3572 4577 3676 4583
rect 3684 4577 3772 4583
rect 3796 4577 3964 4583
rect 4292 4577 4540 4583
rect 4660 4577 4668 4583
rect 4685 4583 4691 4597
rect 4788 4597 5196 4603
rect 5364 4597 5388 4603
rect 5492 4597 5532 4603
rect 5700 4597 5900 4603
rect 6052 4597 7020 4603
rect 7076 4597 7084 4603
rect 7172 4597 7276 4603
rect 4685 4577 4860 4583
rect 4948 4577 5260 4583
rect 5444 4577 5660 4583
rect 5828 4577 6268 4583
rect 6276 4577 6387 4583
rect 2548 4557 2739 4563
rect 2756 4557 2764 4563
rect 2868 4557 3020 4563
rect 3028 4557 3468 4563
rect 3508 4557 3532 4563
rect 3556 4557 3564 4563
rect 3620 4557 3644 4563
rect 3700 4557 3884 4563
rect 3892 4557 4028 4563
rect 4036 4557 4092 4563
rect 4164 4557 4332 4563
rect 4404 4557 4508 4563
rect 4852 4557 4956 4563
rect 5028 4557 5132 4563
rect 5236 4557 5260 4563
rect 5588 4557 5676 4563
rect 5764 4557 6028 4563
rect 6036 4557 6124 4563
rect 6381 4563 6387 4577
rect 6381 4557 6700 4563
rect 148 4537 188 4543
rect 404 4537 476 4543
rect 692 4537 764 4543
rect 1332 4537 1372 4543
rect 1380 4537 1404 4543
rect 1572 4537 1612 4543
rect 1620 4537 1628 4543
rect 1636 4537 1708 4543
rect 2020 4537 2124 4543
rect 2132 4537 2252 4543
rect 2292 4537 2348 4543
rect 2548 4537 2572 4543
rect 2580 4537 2588 4543
rect 2612 4537 2764 4543
rect 2836 4537 2924 4543
rect 3076 4537 3084 4543
rect 3140 4537 3292 4543
rect 3364 4537 3484 4543
rect 3652 4537 4108 4543
rect 4196 4537 4236 4543
rect 4509 4543 4515 4556
rect 4509 4537 5052 4543
rect 5092 4537 5139 4543
rect 5133 4524 5139 4537
rect 5156 4537 5244 4543
rect 5309 4537 5692 4543
rect 5309 4524 5315 4537
rect 5716 4537 5868 4543
rect 5876 4537 5980 4543
rect 6148 4537 6316 4543
rect 6372 4537 6444 4543
rect 6580 4537 6956 4543
rect 6964 4537 7100 4543
rect 20 4517 44 4523
rect 100 4517 204 4523
rect 212 4517 300 4523
rect 852 4517 892 4523
rect 1060 4517 1084 4523
rect 1476 4517 1516 4523
rect 2004 4517 2060 4523
rect 2308 4517 2364 4523
rect 2580 4517 2636 4523
rect 2756 4517 2796 4523
rect 2900 4517 3004 4523
rect 3492 4517 3564 4523
rect 3764 4517 3804 4523
rect 3812 4517 3900 4523
rect 3908 4517 3980 4523
rect 4020 4517 4268 4523
rect 4276 4517 4300 4523
rect 4484 4517 4556 4523
rect 4564 4517 4588 4523
rect 4644 4517 4716 4523
rect 4900 4517 5052 4523
rect 5140 4517 5164 4523
rect 5220 4517 5308 4523
rect 5396 4517 5468 4523
rect 5476 4517 5596 4523
rect 5652 4517 6204 4523
rect 6212 4517 6220 4523
rect 6244 4517 6300 4523
rect 6420 4517 6540 4523
rect 6580 4517 6668 4523
rect 6756 4517 6780 4523
rect 6788 4517 6828 4523
rect 6836 4517 6892 4523
rect 6900 4517 6924 4523
rect 6932 4517 6940 4523
rect 7124 4517 7132 4523
rect 36 4497 92 4503
rect 468 4497 524 4503
rect 964 4497 1132 4503
rect 1140 4497 1180 4503
rect 1556 4497 1692 4503
rect 1908 4497 1932 4503
rect 2052 4497 2716 4503
rect 2724 4497 3004 4503
rect 3012 4497 3036 4503
rect 3060 4497 3356 4503
rect 3460 4497 3468 4503
rect 3540 4497 3596 4503
rect 3764 4497 4060 4503
rect 4708 4497 4796 4503
rect 4820 4497 4892 4503
rect 5124 4497 5292 4503
rect 5364 4497 5804 4503
rect 5908 4497 6044 4503
rect 6068 4497 6284 4503
rect 6324 4497 6636 4503
rect 7156 4497 7212 4503
rect 372 4477 572 4483
rect 1380 4477 1580 4483
rect 1588 4477 1772 4483
rect 1956 4477 2492 4483
rect 3060 4477 3836 4483
rect 3940 4477 3964 4483
rect 4772 4477 4812 4483
rect 4836 4477 4908 4483
rect 5044 4477 5228 4483
rect 5268 4477 6188 4483
rect 6340 4477 6684 4483
rect 1652 4457 1996 4463
rect 2004 4457 2620 4463
rect 2628 4457 3724 4463
rect 3732 4457 3868 4463
rect 3924 4457 3996 4463
rect 5012 4457 5308 4463
rect 5508 4457 5516 4463
rect 5668 4457 6028 4463
rect 6100 4457 6172 4463
rect 6292 4457 6364 4463
rect 6532 4457 6620 4463
rect 6628 4457 7180 4463
rect 1924 4437 2028 4443
rect 2164 4437 2188 4443
rect 2452 4437 2604 4443
rect 2916 4437 3180 4443
rect 3204 4437 3228 4443
rect 3252 4437 3324 4443
rect 3508 4437 4524 4443
rect 4596 4437 5004 4443
rect 5076 4437 5612 4443
rect 6157 4437 6252 4443
rect 6157 4424 6163 4437
rect 1972 4417 2348 4423
rect 2388 4417 3100 4423
rect 3156 4417 3276 4423
rect 4532 4417 5212 4423
rect 5332 4417 5404 4423
rect 5460 4417 5820 4423
rect 5844 4417 6108 4423
rect 6116 4417 6156 4423
rect 6196 4417 6508 4423
rect 1410 4414 1470 4416
rect 1410 4406 1411 4414
rect 1420 4406 1421 4414
rect 1459 4406 1460 4414
rect 1469 4406 1470 4414
rect 1410 4404 1470 4406
rect 4418 4414 4478 4416
rect 4418 4406 4419 4414
rect 4428 4406 4429 4414
rect 4467 4406 4468 4414
rect 4477 4406 4478 4414
rect 4418 4404 4478 4406
rect 516 4397 1148 4403
rect 2084 4397 2252 4403
rect 2564 4397 2700 4403
rect 2708 4397 3420 4403
rect 3444 4397 3500 4403
rect 3796 4397 3948 4403
rect 4772 4397 5020 4403
rect 5060 4397 6316 4403
rect 660 4377 780 4383
rect 788 4377 924 4383
rect 1396 4377 1420 4383
rect 1428 4377 1500 4383
rect 1508 4377 1612 4383
rect 1620 4377 1980 4383
rect 1988 4377 2220 4383
rect 2372 4377 2396 4383
rect 2804 4377 2892 4383
rect 3028 4377 4012 4383
rect 5076 4377 5459 4383
rect 612 4357 748 4363
rect 1332 4357 1436 4363
rect 1444 4357 1660 4363
rect 1668 4357 1868 4363
rect 1988 4357 2044 4363
rect 2180 4357 2236 4363
rect 2356 4357 3084 4363
rect 3092 4357 4028 4363
rect 4116 4357 5436 4363
rect 5453 4363 5459 4377
rect 5812 4377 6092 4383
rect 6132 4377 6156 4383
rect 5453 4357 6236 4363
rect 132 4337 236 4343
rect 276 4337 348 4343
rect 356 4337 620 4343
rect 676 4337 988 4343
rect 1156 4337 1299 4343
rect 1293 4324 1299 4337
rect 1364 4337 1484 4343
rect 1636 4337 1692 4343
rect 1796 4337 1900 4343
rect 2068 4337 2188 4343
rect 2196 4337 3628 4343
rect 3700 4337 4988 4343
rect 5140 4337 5148 4343
rect 5268 4337 5324 4343
rect 5348 4337 5388 4343
rect 5572 4337 5612 4343
rect 5716 4337 6124 4343
rect 6372 4337 6492 4343
rect 6500 4337 6556 4343
rect 148 4317 364 4323
rect 532 4317 556 4323
rect 628 4317 748 4323
rect 884 4317 892 4323
rect 980 4317 1068 4323
rect 1300 4317 2268 4323
rect 2340 4317 2380 4323
rect 2404 4317 2476 4323
rect 2484 4317 2540 4323
rect 2548 4317 2684 4323
rect 2740 4317 2876 4323
rect 3268 4317 3292 4323
rect 3332 4317 3452 4323
rect 3540 4317 3644 4323
rect 4820 4317 5644 4323
rect 5684 4317 5820 4323
rect 5828 4317 6076 4323
rect 6084 4317 6172 4323
rect 6244 4317 6268 4323
rect 6596 4317 6636 4323
rect 6644 4317 6716 4323
rect 6724 4317 6748 4323
rect 6756 4317 6796 4323
rect 6804 4317 6892 4323
rect 7156 4317 7180 4323
rect 292 4297 396 4303
rect 404 4297 700 4303
rect 1060 4297 1068 4303
rect 1076 4297 1180 4303
rect 1188 4297 1228 4303
rect 1268 4297 1372 4303
rect 1540 4297 1580 4303
rect 1748 4297 1932 4303
rect 2132 4297 2140 4303
rect 2212 4297 2236 4303
rect 2404 4297 2428 4303
rect 2580 4297 2604 4303
rect 2612 4297 2652 4303
rect 2900 4297 2988 4303
rect 3396 4297 3436 4303
rect 4164 4297 4188 4303
rect 4804 4297 4844 4303
rect 4852 4297 5036 4303
rect 5092 4297 5484 4303
rect 5492 4297 5548 4303
rect 5588 4297 5612 4303
rect 5652 4297 5756 4303
rect 5876 4297 5884 4303
rect 5892 4297 6252 4303
rect 6500 4297 6588 4303
rect 6788 4297 7052 4303
rect 7188 4297 7308 4303
rect 116 4277 172 4283
rect 500 4277 604 4283
rect 660 4277 748 4283
rect 756 4277 908 4283
rect 916 4277 924 4283
rect 1220 4277 1324 4283
rect 1380 4277 1708 4283
rect 1732 4277 1772 4283
rect 1828 4277 1884 4283
rect 1924 4277 2204 4283
rect 2212 4277 2364 4283
rect 2468 4277 2508 4283
rect 2653 4277 2780 4283
rect 52 4257 140 4263
rect 228 4257 316 4263
rect 324 4257 380 4263
rect 436 4257 508 4263
rect 612 4257 1180 4263
rect 1188 4257 1308 4263
rect 1316 4257 1740 4263
rect 1828 4257 1868 4263
rect 1876 4257 2012 4263
rect 2164 4257 2316 4263
rect 2653 4263 2659 4277
rect 3348 4277 3404 4283
rect 3428 4277 3596 4283
rect 3709 4283 3715 4296
rect 3709 4277 3724 4283
rect 4244 4277 4332 4283
rect 4340 4277 4444 4283
rect 4452 4277 4652 4283
rect 4884 4277 4892 4283
rect 4964 4277 5116 4283
rect 5316 4277 5340 4283
rect 5540 4277 5708 4283
rect 5748 4277 5884 4283
rect 5892 4277 5916 4283
rect 5924 4277 6332 4283
rect 6340 4277 6492 4283
rect 6580 4277 6620 4283
rect 6628 4277 6652 4283
rect 6820 4277 6844 4283
rect 6964 4277 7132 4283
rect 7156 4277 7180 4283
rect 2356 4257 2659 4263
rect 2676 4257 2748 4263
rect 3188 4257 3708 4263
rect 3716 4257 3724 4263
rect 3972 4257 4156 4263
rect 4164 4257 4316 4263
rect 5028 4257 5132 4263
rect 5204 4257 5324 4263
rect 5348 4257 5356 4263
rect 5428 4257 5564 4263
rect 5604 4257 5644 4263
rect 5732 4257 5740 4263
rect 5876 4257 6044 4263
rect 6228 4257 6300 4263
rect 6532 4257 6652 4263
rect 372 4237 412 4243
rect 420 4237 620 4243
rect 676 4237 860 4243
rect 900 4237 1004 4243
rect 1140 4237 1196 4243
rect 1716 4237 1756 4243
rect 1780 4237 1836 4243
rect 2260 4237 2428 4243
rect 2468 4237 2524 4243
rect 2532 4237 2588 4243
rect 2996 4237 3340 4243
rect 3508 4237 3532 4243
rect 4580 4237 4604 4243
rect 4612 4237 4636 4243
rect 4644 4237 4780 4243
rect 5300 4237 5372 4243
rect 5508 4237 5548 4243
rect 5620 4237 5644 4243
rect 5732 4237 5852 4243
rect 6228 4237 6716 4243
rect 6724 4237 6940 4243
rect 788 4217 1052 4223
rect 1236 4217 1276 4223
rect 1412 4217 1644 4223
rect 2420 4217 2476 4223
rect 2484 4217 2780 4223
rect 3092 4217 3100 4223
rect 3236 4217 3516 4223
rect 3748 4217 4092 4223
rect 5476 4217 5852 4223
rect 6020 4217 6220 4223
rect 6356 4217 6444 4223
rect 6452 4217 6924 4223
rect 2914 4214 2974 4216
rect 2914 4206 2915 4214
rect 2924 4206 2925 4214
rect 2963 4206 2964 4214
rect 2973 4206 2974 4214
rect 2914 4204 2974 4206
rect 5922 4214 5982 4216
rect 5922 4206 5923 4214
rect 5932 4206 5933 4214
rect 5971 4206 5972 4214
rect 5981 4206 5982 4214
rect 5922 4204 5982 4206
rect 68 4197 236 4203
rect 244 4197 460 4203
rect 708 4197 972 4203
rect 996 4197 1116 4203
rect 1444 4197 1964 4203
rect 2228 4197 2252 4203
rect 2580 4197 2732 4203
rect 3380 4197 3404 4203
rect 3636 4197 4028 4203
rect 4596 4197 4732 4203
rect 4740 4197 4780 4203
rect 5012 4197 5148 4203
rect 5156 4197 5356 4203
rect 5396 4197 5532 4203
rect 5540 4197 5580 4203
rect 5620 4197 5740 4203
rect 5764 4197 5836 4203
rect 6212 4197 6300 4203
rect 6308 4197 6508 4203
rect 6580 4197 6828 4203
rect 116 4177 460 4183
rect 708 4177 1004 4183
rect 1012 4177 1020 4183
rect 1060 4177 1948 4183
rect 2228 4177 2252 4183
rect 2276 4177 2476 4183
rect 2708 4177 2764 4183
rect 2804 4177 2908 4183
rect 2916 4177 3740 4183
rect 3796 4177 3820 4183
rect 3988 4177 4076 4183
rect 4724 4177 4828 4183
rect 4932 4177 5132 4183
rect 5140 4177 5180 4183
rect 5572 4177 6028 4183
rect 6036 4177 6284 4183
rect 6324 4177 6348 4183
rect 6372 4177 6908 4183
rect 6932 4177 6972 4183
rect 164 4157 540 4163
rect 836 4157 924 4163
rect 948 4157 1308 4163
rect 1716 4157 1820 4163
rect 1828 4157 1980 4163
rect 1988 4157 2108 4163
rect 2244 4157 2460 4163
rect 2532 4157 2620 4163
rect 2836 4157 2860 4163
rect 2868 4157 2924 4163
rect 3709 4157 4108 4163
rect 3709 4144 3715 4157
rect 4116 4157 4188 4163
rect 4484 4157 4684 4163
rect 4692 4157 4876 4163
rect 4900 4157 4972 4163
rect 5236 4157 5276 4163
rect 5300 4157 5612 4163
rect 5668 4157 5772 4163
rect 5780 4157 5836 4163
rect 5892 4157 5932 4163
rect 6084 4157 6156 4163
rect 6276 4157 6812 4163
rect 532 4137 732 4143
rect 788 4137 812 4143
rect 964 4137 1084 4143
rect 1092 4137 1164 4143
rect 1188 4137 1436 4143
rect 1604 4137 1900 4143
rect 1908 4137 2188 4143
rect 2196 4137 2316 4143
rect 2436 4137 2556 4143
rect 2580 4137 2636 4143
rect 2788 4137 2828 4143
rect 3300 4137 3388 4143
rect 3396 4137 3404 4143
rect 3476 4137 3500 4143
rect 3508 4137 3548 4143
rect 3556 4137 3612 4143
rect 3620 4137 3692 4143
rect 3700 4137 3708 4143
rect 3892 4137 3948 4143
rect 4372 4137 4396 4143
rect 4756 4137 5020 4143
rect 5236 4137 5388 4143
rect 5396 4137 5644 4143
rect 5652 4137 5724 4143
rect 5780 4137 5884 4143
rect 5892 4137 6284 4143
rect 6324 4137 6412 4143
rect 6756 4137 7052 4143
rect 52 4117 76 4123
rect 852 4117 972 4123
rect 1028 4117 1084 4123
rect 1284 4117 1340 4123
rect 1588 4117 1692 4123
rect 2132 4117 2236 4123
rect 2244 4117 2284 4123
rect 2292 4117 2348 4123
rect 2420 4117 2540 4123
rect 2660 4117 2748 4123
rect 2756 4117 2812 4123
rect 3044 4117 3244 4123
rect 3252 4117 3484 4123
rect 3620 4117 3628 4123
rect 3684 4117 3740 4123
rect 3876 4117 3884 4123
rect 3892 4117 4140 4123
rect 4500 4117 4540 4123
rect 4612 4117 4876 4123
rect 4884 4117 4988 4123
rect 5620 4117 5868 4123
rect 5892 4117 5948 4123
rect 6052 4117 6092 4123
rect 6132 4117 6172 4123
rect 6260 4117 6540 4123
rect 6884 4117 7084 4123
rect 7252 4117 7260 4123
rect 148 4097 220 4103
rect 1060 4097 1068 4103
rect 1172 4097 1660 4103
rect 1748 4097 1852 4103
rect 1988 4097 2284 4103
rect 2292 4097 2988 4103
rect 3092 4097 3148 4103
rect 3236 4097 3244 4103
rect 3869 4103 3875 4116
rect 3508 4097 3875 4103
rect 4212 4097 4780 4103
rect 4820 4097 4860 4103
rect 4964 4097 5052 4103
rect 5252 4097 5308 4103
rect 5396 4097 5452 4103
rect 5460 4097 5676 4103
rect 5700 4097 5804 4103
rect 5812 4097 6476 4103
rect 6564 4097 6700 4103
rect 6804 4097 6940 4103
rect 7044 4097 7084 4103
rect 36 4077 92 4083
rect 1012 4077 1132 4083
rect 1140 4077 1580 4083
rect 2388 4077 2412 4083
rect 2484 4077 2572 4083
rect 2852 4077 3036 4083
rect 3076 4077 3084 4083
rect 3444 4077 3820 4083
rect 4020 4077 4124 4083
rect 4868 4077 4908 4083
rect 4948 4077 5292 4083
rect 5412 4077 5660 4083
rect 5716 4077 5788 4083
rect 5844 4077 6028 4083
rect 6052 4077 6300 4083
rect 6516 4077 6588 4083
rect 6660 4077 6780 4083
rect 6948 4077 7164 4083
rect 916 4057 1276 4063
rect 1332 4057 1516 4063
rect 2036 4057 2060 4063
rect 2612 4057 3052 4063
rect 3060 4057 3116 4063
rect 3572 4057 4908 4063
rect 5524 4057 5612 4063
rect 5629 4057 6092 4063
rect 212 4037 236 4043
rect 612 4037 876 4043
rect 884 4037 1132 4043
rect 1140 4037 2044 4043
rect 2740 4037 3324 4043
rect 3332 4037 3756 4043
rect 3764 4037 4012 4043
rect 5629 4043 5635 4057
rect 6196 4057 6252 4063
rect 6260 4057 6428 4063
rect 6436 4057 6444 4063
rect 7140 4057 7148 4063
rect 5268 4037 5635 4043
rect 5796 4037 6460 4043
rect 6468 4037 6924 4043
rect 436 4017 636 4023
rect 644 4017 908 4023
rect 916 4017 1148 4023
rect 1492 4017 2028 4023
rect 2676 4017 2732 4023
rect 2740 4017 2876 4023
rect 3156 4017 3676 4023
rect 4516 4017 6044 4023
rect 6068 4017 6268 4023
rect 6276 4017 6316 4023
rect 6900 4017 7196 4023
rect 7220 4017 7276 4023
rect 1410 4014 1470 4016
rect 1410 4006 1411 4014
rect 1420 4006 1421 4014
rect 1459 4006 1460 4014
rect 1469 4006 1470 4014
rect 1410 4004 1470 4006
rect 4418 4014 4478 4016
rect 4418 4006 4419 4014
rect 4428 4006 4429 4014
rect 4467 4006 4468 4014
rect 4477 4006 4478 4014
rect 4418 4004 4478 4006
rect 868 3997 1100 4003
rect 1172 3997 1388 4003
rect 2516 3997 2732 4003
rect 2740 3997 2844 4003
rect 3044 3997 3452 4003
rect 3476 3997 4220 4003
rect 4228 3997 4284 4003
rect 4532 3997 6044 4003
rect 6132 3997 6220 4003
rect 6260 3997 6396 4003
rect 6484 3997 6700 4003
rect 1364 3977 1644 3983
rect 1892 3977 3139 3983
rect 900 3957 2108 3963
rect 2996 3957 3084 3963
rect 3133 3963 3139 3977
rect 3156 3977 3212 3983
rect 3316 3977 3436 3983
rect 3476 3977 3532 3983
rect 3604 3977 3820 3983
rect 4100 3977 4188 3983
rect 4596 3977 4652 3983
rect 4660 3977 4732 3983
rect 4740 3977 5244 3983
rect 5540 3977 5724 3983
rect 5796 3977 5916 3983
rect 5924 3977 6620 3983
rect 3133 3957 3196 3963
rect 3220 3957 3276 3963
rect 3284 3957 3468 3963
rect 3732 3957 4508 3963
rect 5684 3957 6028 3963
rect 6052 3957 6156 3963
rect 6196 3957 6243 3963
rect 20 3937 44 3943
rect 628 3937 684 3943
rect 692 3937 860 3943
rect 868 3937 1180 3943
rect 1364 3937 1372 3943
rect 1476 3937 1532 3943
rect 1684 3937 1996 3943
rect 2068 3937 2284 3943
rect 2292 3937 2364 3943
rect 2372 3937 2508 3943
rect 4948 3937 5116 3943
rect 5133 3937 5260 3943
rect 52 3917 124 3923
rect 180 3917 252 3923
rect 356 3917 540 3923
rect 548 3917 572 3923
rect 660 3917 700 3923
rect 788 3917 812 3923
rect 1300 3917 1555 3923
rect 1549 3904 1555 3917
rect 1716 3917 1820 3923
rect 1828 3917 1948 3923
rect 2004 3917 2620 3923
rect 2804 3917 3036 3923
rect 3924 3917 4108 3923
rect 4180 3917 4252 3923
rect 4916 3917 4988 3923
rect 5133 3923 5139 3937
rect 5300 3937 5484 3943
rect 5668 3937 5772 3943
rect 6116 3937 6220 3943
rect 6237 3943 6243 3957
rect 6276 3957 6684 3963
rect 6237 3937 6380 3943
rect 6420 3937 6508 3943
rect 6580 3937 6748 3943
rect 6756 3937 6860 3943
rect 5028 3917 5139 3923
rect 5220 3917 5324 3923
rect 5604 3917 5772 3923
rect 5892 3917 6060 3923
rect 6148 3917 6252 3923
rect 6292 3917 6364 3923
rect 6372 3917 6444 3923
rect 6461 3917 6508 3923
rect 68 3897 124 3903
rect 132 3897 156 3903
rect 244 3897 460 3903
rect 484 3897 764 3903
rect 916 3897 924 3903
rect 1124 3897 1196 3903
rect 1204 3897 1260 3903
rect 1284 3897 1388 3903
rect 1572 3897 1676 3903
rect 1700 3897 1900 3903
rect 1940 3897 1980 3903
rect 2020 3897 2188 3903
rect 2196 3897 2236 3903
rect 2564 3897 2572 3903
rect 2708 3897 2844 3903
rect 3044 3897 3132 3903
rect 3140 3897 3180 3903
rect 3604 3897 3660 3903
rect 4420 3897 4444 3903
rect 4676 3897 4700 3903
rect 4964 3897 5084 3903
rect 5108 3897 5196 3903
rect 5204 3897 5500 3903
rect 5508 3897 5836 3903
rect 6461 3903 6467 3917
rect 6548 3917 6812 3923
rect 6836 3917 6972 3923
rect 7156 3917 7180 3923
rect 5988 3897 6467 3903
rect 6500 3897 6652 3903
rect 6788 3897 6828 3903
rect 6900 3897 7100 3903
rect 7156 3897 7196 3903
rect 7236 3897 7276 3903
rect 116 3877 236 3883
rect 292 3877 364 3883
rect 532 3877 716 3883
rect 852 3877 1731 3883
rect 1069 3864 1075 3877
rect 1725 3864 1731 3877
rect 2324 3877 2380 3883
rect 2388 3877 2604 3883
rect 2612 3877 2636 3883
rect 2644 3877 2652 3883
rect 2724 3877 2764 3883
rect 2772 3877 2860 3883
rect 2884 3877 3004 3883
rect 3012 3877 3052 3883
rect 3332 3877 3436 3883
rect 3812 3877 3868 3883
rect 3892 3877 4028 3883
rect 4052 3877 4156 3883
rect 4868 3877 5324 3883
rect 5428 3877 5532 3883
rect 5780 3877 5820 3883
rect 5956 3877 6268 3883
rect 6484 3877 6492 3883
rect 6628 3877 6668 3883
rect 6676 3877 6892 3883
rect 7028 3877 7260 3883
rect 276 3857 300 3863
rect 308 3857 460 3863
rect 468 3857 540 3863
rect 580 3857 652 3863
rect 724 3857 876 3863
rect 980 3857 1020 3863
rect 1245 3857 1564 3863
rect 196 3837 220 3843
rect 340 3837 860 3843
rect 1245 3843 1251 3857
rect 1732 3857 1836 3863
rect 2148 3857 2284 3863
rect 2996 3857 3164 3863
rect 3268 3857 3292 3863
rect 3300 3857 3324 3863
rect 3748 3857 3932 3863
rect 3940 3857 4076 3863
rect 4852 3857 4956 3863
rect 4980 3857 5036 3863
rect 5044 3857 5228 3863
rect 5284 3857 5420 3863
rect 5460 3857 5692 3863
rect 5764 3857 5804 3863
rect 5812 3857 6108 3863
rect 6244 3857 6252 3863
rect 6308 3857 6492 3863
rect 6548 3857 6700 3863
rect 6948 3857 7052 3863
rect 7092 3857 7292 3863
rect 1012 3837 1251 3843
rect 1268 3837 1324 3843
rect 2461 3837 2620 3843
rect 2461 3824 2467 3837
rect 3012 3837 3148 3843
rect 3236 3837 3260 3843
rect 3268 3837 3564 3843
rect 3796 3837 3884 3843
rect 4212 3837 4476 3843
rect 4548 3837 4764 3843
rect 4772 3837 5212 3843
rect 5252 3837 5484 3843
rect 5700 3837 5884 3843
rect 6068 3837 6444 3843
rect 6452 3837 6620 3843
rect 6628 3837 6636 3843
rect 6644 3837 6732 3843
rect 6740 3837 6956 3843
rect 7252 3837 7260 3843
rect 196 3817 316 3823
rect 740 3817 764 3823
rect 772 3817 812 3823
rect 820 3817 828 3823
rect 836 3817 972 3823
rect 980 3817 1692 3823
rect 2052 3817 2460 3823
rect 2477 3817 2780 3823
rect 820 3797 908 3803
rect 1300 3797 1468 3803
rect 1956 3797 1996 3803
rect 2004 3797 2204 3803
rect 2228 3797 2268 3803
rect 2477 3803 2483 3817
rect 4900 3817 4908 3823
rect 4980 3817 5084 3823
rect 5092 3817 5180 3823
rect 5236 3817 5260 3823
rect 5284 3817 5340 3823
rect 5524 3817 5564 3823
rect 5572 3817 5756 3823
rect 6020 3817 6076 3823
rect 6084 3817 6412 3823
rect 6420 3817 6556 3823
rect 6948 3817 6956 3823
rect 7044 3817 7084 3823
rect 2914 3814 2974 3816
rect 2914 3806 2915 3814
rect 2924 3806 2925 3814
rect 2963 3806 2964 3814
rect 2973 3806 2974 3814
rect 2914 3804 2974 3806
rect 5922 3814 5982 3816
rect 5922 3806 5923 3814
rect 5932 3806 5933 3814
rect 5971 3806 5972 3814
rect 5981 3806 5982 3814
rect 5922 3804 5982 3806
rect 2324 3797 2483 3803
rect 2516 3797 2668 3803
rect 2788 3797 2876 3803
rect 3588 3797 3596 3803
rect 3860 3797 3900 3803
rect 4132 3797 4204 3803
rect 4244 3797 4268 3803
rect 4308 3797 4348 3803
rect 4420 3797 4604 3803
rect 4708 3797 4748 3803
rect 4804 3797 5068 3803
rect 5092 3797 5116 3803
rect 5172 3797 5420 3803
rect 6068 3797 6140 3803
rect 6180 3797 6572 3803
rect 6996 3797 7084 3803
rect 436 3777 476 3783
rect 996 3777 1027 3783
rect 68 3757 252 3763
rect 468 3757 524 3763
rect 564 3757 716 3763
rect 788 3757 844 3763
rect 884 3757 940 3763
rect 1021 3763 1027 3777
rect 1108 3777 1676 3783
rect 1732 3777 2268 3783
rect 2644 3777 3052 3783
rect 3108 3777 3212 3783
rect 3396 3777 3500 3783
rect 3524 3777 3596 3783
rect 3604 3777 3724 3783
rect 3732 3777 3772 3783
rect 3844 3777 3852 3783
rect 4100 3777 4220 3783
rect 4308 3777 4588 3783
rect 4900 3777 4972 3783
rect 5028 3777 5596 3783
rect 5604 3777 5612 3783
rect 5652 3777 5756 3783
rect 5901 3783 5907 3796
rect 5901 3777 5948 3783
rect 5972 3777 6028 3783
rect 6116 3777 6156 3783
rect 6260 3777 6348 3783
rect 6484 3777 6716 3783
rect 6733 3777 6908 3783
rect 1021 3757 1324 3763
rect 1844 3757 1980 3763
rect 2260 3757 2355 3763
rect 244 3737 284 3743
rect 292 3737 396 3743
rect 420 3737 476 3743
rect 564 3737 915 3743
rect 909 3724 915 3737
rect 1188 3737 1244 3743
rect 1348 3737 1356 3743
rect 1924 3737 2012 3743
rect 2148 3737 2204 3743
rect 2324 3737 2332 3743
rect 2349 3743 2355 3757
rect 2452 3757 2876 3763
rect 3364 3757 3676 3763
rect 3684 3757 3692 3763
rect 3764 3757 3804 3763
rect 3828 3757 3852 3763
rect 4068 3757 4108 3763
rect 4116 3757 4172 3763
rect 4180 3757 4236 3763
rect 4276 3757 4524 3763
rect 5060 3757 5148 3763
rect 5204 3757 5276 3763
rect 5332 3757 6252 3763
rect 6733 3763 6739 3777
rect 7076 3777 7340 3783
rect 6388 3757 6739 3763
rect 6852 3757 7004 3763
rect 7188 3757 7228 3763
rect 7252 3757 7340 3763
rect 2349 3737 2412 3743
rect 2564 3737 2716 3743
rect 2756 3737 2812 3743
rect 2916 3737 3036 3743
rect 3236 3737 3340 3743
rect 3508 3737 3708 3743
rect 3716 3737 3996 3743
rect 4004 3737 4252 3743
rect 4260 3737 4332 3743
rect 4356 3737 4412 3743
rect 4580 3737 4636 3743
rect 4676 3737 4700 3743
rect 4788 3737 4940 3743
rect 5044 3737 5164 3743
rect 5172 3737 5196 3743
rect 5332 3737 5388 3743
rect 5428 3737 5468 3743
rect 5476 3737 5644 3743
rect 5748 3737 5868 3743
rect 6068 3737 6092 3743
rect 6404 3737 6476 3743
rect 6484 3737 6652 3743
rect 6660 3737 6844 3743
rect 6932 3737 7052 3743
rect 7092 3737 7196 3743
rect 116 3717 156 3723
rect 164 3717 172 3723
rect 516 3717 604 3723
rect 660 3717 668 3723
rect 820 3717 844 3723
rect 916 3717 1724 3723
rect 1828 3717 1884 3723
rect 2004 3717 2156 3723
rect 2308 3717 2348 3723
rect 2484 3717 2492 3723
rect 2532 3717 2604 3723
rect 2628 3717 2636 3723
rect 3316 3717 3340 3723
rect 3364 3717 3404 3723
rect 3460 3717 3692 3723
rect 3748 3717 3820 3723
rect 3876 3717 3932 3723
rect 3940 3717 3980 3723
rect 4036 3717 4268 3723
rect 4292 3717 4588 3723
rect 4932 3717 4940 3723
rect 5012 3717 5036 3723
rect 5108 3717 5180 3723
rect 5252 3717 5452 3723
rect 5508 3717 5532 3723
rect 5684 3717 5724 3723
rect 5805 3717 6044 3723
rect 404 3697 428 3703
rect 596 3697 876 3703
rect 1236 3697 1276 3703
rect 1380 3697 1500 3703
rect 1508 3697 1564 3703
rect 1572 3697 1644 3703
rect 1821 3703 1827 3716
rect 1652 3697 1827 3703
rect 1908 3697 2124 3703
rect 3044 3697 3340 3703
rect 3428 3697 3539 3703
rect 589 3683 595 3696
rect 324 3677 595 3683
rect 836 3677 972 3683
rect 1396 3677 1628 3683
rect 1668 3677 3068 3683
rect 3188 3677 3436 3683
rect 3460 3677 3516 3683
rect 3533 3683 3539 3697
rect 3556 3697 3756 3703
rect 4052 3697 4300 3703
rect 4308 3697 4380 3703
rect 5108 3697 5116 3703
rect 5284 3697 5404 3703
rect 5412 3697 5420 3703
rect 5805 3703 5811 3717
rect 6052 3717 6188 3723
rect 6324 3717 6588 3723
rect 6596 3717 6668 3723
rect 6724 3717 6796 3723
rect 6820 3717 6956 3723
rect 6964 3717 7132 3723
rect 7284 3717 7324 3723
rect 7332 3717 7372 3723
rect 5524 3697 5811 3703
rect 5844 3697 6012 3703
rect 6036 3697 6428 3703
rect 6436 3697 6444 3703
rect 6548 3697 6620 3703
rect 6660 3697 6764 3703
rect 6884 3697 6972 3703
rect 7277 3703 7283 3716
rect 6996 3697 7283 3703
rect 3533 3677 3580 3683
rect 3972 3677 4108 3683
rect 4116 3677 4124 3683
rect 4148 3677 4396 3683
rect 4612 3677 4732 3683
rect 4916 3677 5356 3683
rect 5636 3677 5836 3683
rect 5844 3677 6076 3683
rect 6164 3677 6300 3683
rect 6356 3677 6604 3683
rect 6708 3677 6732 3683
rect 6740 3677 7100 3683
rect 532 3657 1260 3663
rect 1396 3657 1516 3663
rect 1524 3657 1580 3663
rect 2116 3657 2204 3663
rect 2212 3657 2364 3663
rect 2372 3657 2396 3663
rect 3332 3657 3740 3663
rect 3748 3657 3948 3663
rect 4388 3657 4444 3663
rect 4996 3657 5084 3663
rect 5108 3657 5292 3663
rect 5652 3657 6028 3663
rect 6052 3657 6076 3663
rect 6100 3657 6220 3663
rect 6340 3657 6796 3663
rect 6932 3657 7020 3663
rect 7076 3657 7164 3663
rect 596 3637 620 3643
rect 852 3637 1356 3643
rect 1476 3637 1596 3643
rect 2644 3637 2668 3643
rect 3604 3637 3612 3643
rect 3709 3637 4220 3643
rect 820 3617 1052 3623
rect 1588 3617 1740 3623
rect 3709 3623 3715 3637
rect 4884 3637 5580 3643
rect 5748 3637 6188 3643
rect 6212 3637 6220 3643
rect 6708 3637 6764 3643
rect 6916 3637 7116 3643
rect 3492 3617 3715 3623
rect 3732 3617 3868 3623
rect 4772 3617 4812 3623
rect 4820 3617 6716 3623
rect 6724 3617 6780 3623
rect 6836 3617 6988 3623
rect 7012 3617 7116 3623
rect 1410 3614 1470 3616
rect 1410 3606 1411 3614
rect 1420 3606 1421 3614
rect 1459 3606 1460 3614
rect 1469 3606 1470 3614
rect 1410 3604 1470 3606
rect 4418 3614 4478 3616
rect 4418 3606 4419 3614
rect 4428 3606 4429 3614
rect 4467 3606 4468 3614
rect 4477 3606 4478 3614
rect 4418 3604 4478 3606
rect 692 3597 732 3603
rect 1652 3597 1676 3603
rect 3380 3597 3436 3603
rect 3540 3597 4300 3603
rect 5684 3597 5980 3603
rect 6020 3597 6492 3603
rect 6772 3597 7052 3603
rect 68 3577 172 3583
rect 180 3577 284 3583
rect 292 3577 556 3583
rect 1332 3577 1443 3583
rect 756 3557 796 3563
rect 948 3557 1020 3563
rect 1124 3557 1276 3563
rect 1380 3557 1404 3563
rect 1437 3563 1443 3577
rect 1460 3577 1628 3583
rect 1636 3577 1804 3583
rect 1812 3577 1868 3583
rect 1892 3577 1932 3583
rect 3444 3577 3484 3583
rect 3764 3577 3980 3583
rect 4484 3577 4652 3583
rect 5588 3577 6572 3583
rect 6580 3577 7052 3583
rect 7060 3577 7180 3583
rect 1437 3557 1900 3563
rect 2308 3557 2524 3563
rect 2852 3557 2883 3563
rect 308 3537 332 3543
rect 340 3537 412 3543
rect 420 3537 460 3543
rect 516 3537 1180 3543
rect 1236 3537 1372 3543
rect 1556 3537 1580 3543
rect 1780 3537 1804 3543
rect 2260 3537 2364 3543
rect 2580 3537 2732 3543
rect 2740 3537 2860 3543
rect 2877 3543 2883 3557
rect 3732 3557 3820 3563
rect 3940 3557 3996 3563
rect 4420 3557 4572 3563
rect 5428 3557 5692 3563
rect 5716 3557 5811 3563
rect 2877 3537 3948 3543
rect 3956 3537 3996 3543
rect 4020 3537 4076 3543
rect 4132 3537 4172 3543
rect 4676 3537 4812 3543
rect 5588 3537 5788 3543
rect 5805 3543 5811 3557
rect 6036 3557 6060 3563
rect 6100 3557 6348 3563
rect 6404 3557 6668 3563
rect 6884 3557 6924 3563
rect 7028 3557 7212 3563
rect 5805 3537 6364 3543
rect 6372 3537 6636 3543
rect 6644 3537 6684 3543
rect 6900 3537 6924 3543
rect 6932 3537 7180 3543
rect 756 3517 1084 3523
rect 1172 3517 1196 3523
rect 1524 3517 1548 3523
rect 1620 3517 1628 3523
rect 1636 3517 1884 3523
rect 2052 3517 2076 3523
rect 2308 3517 2460 3523
rect 2484 3517 2492 3523
rect 3108 3517 3292 3523
rect 3460 3517 3596 3523
rect 3604 3517 3788 3523
rect 3796 3517 3852 3523
rect 3860 3517 4092 3523
rect 4100 3517 4108 3523
rect 4772 3517 4812 3523
rect 6068 3517 6188 3523
rect 6196 3517 6220 3523
rect 6548 3517 6652 3523
rect 6868 3517 7020 3523
rect 7140 3517 7372 3523
rect 100 3497 220 3503
rect 228 3497 252 3503
rect 260 3497 316 3503
rect 708 3497 716 3503
rect 724 3497 812 3503
rect 900 3497 924 3503
rect 980 3497 1004 3503
rect 1172 3497 1260 3503
rect 1300 3497 1388 3503
rect 1492 3497 1516 3503
rect 1732 3497 1948 3503
rect 2068 3497 2076 3503
rect 2084 3497 2236 3503
rect 2244 3497 2332 3503
rect 2340 3497 2364 3503
rect 2564 3497 2588 3503
rect 2692 3497 2700 3503
rect 3476 3497 3788 3503
rect 3844 3497 3916 3503
rect 3988 3497 4044 3503
rect 4116 3497 4172 3503
rect 4180 3497 4220 3503
rect 4308 3497 4396 3503
rect 4404 3497 4620 3503
rect 4660 3497 4828 3503
rect 4852 3497 5116 3503
rect 5124 3497 5228 3503
rect 5268 3497 5292 3503
rect 5444 3497 5516 3503
rect 5524 3497 5708 3503
rect 5716 3497 5756 3503
rect 5796 3497 5820 3503
rect 5828 3497 5996 3503
rect 6004 3497 6028 3503
rect 6052 3497 6060 3503
rect 6116 3497 6220 3503
rect 6420 3497 6476 3503
rect 6484 3497 6604 3503
rect 6756 3497 6892 3503
rect 7172 3497 7292 3503
rect 36 3477 108 3483
rect 308 3477 332 3483
rect 340 3477 428 3483
rect 580 3477 764 3483
rect 893 3483 899 3496
rect 772 3477 899 3483
rect 948 3477 1052 3483
rect 1284 3477 1340 3483
rect 1348 3477 1388 3483
rect 1949 3483 1955 3496
rect 1949 3477 1964 3483
rect 2324 3477 2332 3483
rect 2500 3477 2508 3483
rect 2580 3477 2732 3483
rect 2852 3477 3020 3483
rect 3156 3477 3244 3483
rect 3252 3477 3356 3483
rect 3412 3477 3468 3483
rect 3476 3477 3516 3483
rect 3604 3477 3676 3483
rect 3716 3477 3884 3483
rect 3908 3477 4044 3483
rect 4740 3477 4924 3483
rect 5108 3477 5132 3483
rect 5140 3477 5388 3483
rect 5396 3477 5484 3483
rect 5540 3477 5612 3483
rect 5652 3477 5804 3483
rect 5812 3477 6028 3483
rect 6820 3477 6892 3483
rect 6900 3477 7132 3483
rect 7140 3477 7244 3483
rect 180 3457 204 3463
rect 564 3457 748 3463
rect 756 3457 860 3463
rect 868 3457 908 3463
rect 964 3457 1116 3463
rect 1220 3457 1340 3463
rect 1357 3457 1756 3463
rect 884 3437 972 3443
rect 1357 3443 1363 3457
rect 1956 3457 2220 3463
rect 2356 3457 2508 3463
rect 3380 3457 3388 3463
rect 3396 3457 3404 3463
rect 3428 3457 3484 3463
rect 3556 3457 3740 3463
rect 3748 3457 3836 3463
rect 3860 3457 3932 3463
rect 3956 3457 4284 3463
rect 4292 3457 4604 3463
rect 5028 3457 5164 3463
rect 5172 3457 5404 3463
rect 5412 3457 5452 3463
rect 5645 3463 5651 3476
rect 5460 3457 5651 3463
rect 5972 3457 6108 3463
rect 6132 3457 6220 3463
rect 6852 3457 6876 3463
rect 7012 3457 7036 3463
rect 1300 3437 1363 3443
rect 1716 3437 2188 3443
rect 2196 3437 2300 3443
rect 3076 3437 3452 3443
rect 3652 3437 3740 3443
rect 4548 3437 4732 3443
rect 4932 3437 5628 3443
rect 5636 3437 5692 3443
rect 5700 3437 6156 3443
rect 6164 3437 6700 3443
rect 6708 3437 6908 3443
rect 6916 3437 7036 3443
rect 180 3417 2012 3423
rect 2244 3417 2476 3423
rect 3140 3417 3276 3423
rect 3284 3417 3500 3423
rect 4500 3417 4540 3423
rect 4628 3417 4684 3423
rect 5300 3417 5452 3423
rect 5572 3417 5900 3423
rect 6036 3417 6252 3423
rect 6484 3417 7116 3423
rect 2914 3414 2974 3416
rect 2914 3406 2915 3414
rect 2924 3406 2925 3414
rect 2963 3406 2964 3414
rect 2973 3406 2974 3414
rect 2914 3404 2974 3406
rect 5922 3414 5982 3416
rect 5922 3406 5923 3414
rect 5932 3406 5933 3414
rect 5971 3406 5972 3414
rect 5981 3406 5982 3414
rect 5922 3404 5982 3406
rect 500 3397 652 3403
rect 788 3397 812 3403
rect 884 3397 1708 3403
rect 1716 3397 1900 3403
rect 1908 3397 1916 3403
rect 3684 3397 3932 3403
rect 4532 3397 4556 3403
rect 4836 3397 4908 3403
rect 4916 3397 4972 3403
rect 4980 3397 5180 3403
rect 5188 3397 5420 3403
rect 6100 3397 6188 3403
rect 6324 3397 6444 3403
rect 500 3377 924 3383
rect 941 3377 1212 3383
rect 292 3357 524 3363
rect 564 3357 620 3363
rect 788 3357 796 3363
rect 941 3363 947 3377
rect 1636 3377 1708 3383
rect 1828 3377 1884 3383
rect 2084 3377 2460 3383
rect 2868 3377 2972 3383
rect 3396 3377 3900 3383
rect 4020 3377 4284 3383
rect 4580 3377 4764 3383
rect 4772 3377 4860 3383
rect 4868 3377 5004 3383
rect 5044 3377 5084 3383
rect 5092 3377 5340 3383
rect 5348 3377 5372 3383
rect 5732 3377 6092 3383
rect 6132 3377 6492 3383
rect 6772 3377 6844 3383
rect 7140 3377 7212 3383
rect 852 3357 947 3363
rect 1076 3357 1228 3363
rect 1316 3357 1484 3363
rect 1604 3357 1932 3363
rect 2196 3357 2252 3363
rect 2580 3357 2620 3363
rect 2708 3357 2716 3363
rect 2948 3357 3116 3363
rect 3124 3357 3196 3363
rect 3300 3357 3340 3363
rect 3348 3357 3532 3363
rect 3556 3357 3644 3363
rect 3700 3357 3708 3363
rect 3716 3357 3724 3363
rect 3972 3357 4060 3363
rect 4244 3357 4364 3363
rect 4964 3357 5068 3363
rect 5076 3357 5100 3363
rect 5156 3357 5452 3363
rect 5604 3357 5788 3363
rect 6196 3357 6380 3363
rect 7172 3357 7212 3363
rect 52 3337 124 3343
rect 276 3337 332 3343
rect 436 3337 1020 3343
rect 1220 3337 1356 3343
rect 1508 3337 1820 3343
rect 2020 3337 2236 3343
rect 2404 3337 2428 3343
rect 2644 3337 2684 3343
rect 3524 3337 3564 3343
rect 4052 3337 4108 3343
rect 4260 3337 4348 3343
rect 4356 3337 4412 3343
rect 4516 3337 4636 3343
rect 4708 3337 4796 3343
rect 4804 3337 5212 3343
rect 5220 3337 5404 3343
rect 5412 3337 5756 3343
rect 6132 3337 6412 3343
rect 6420 3337 6460 3343
rect 6548 3337 6988 3343
rect 7172 3337 7292 3343
rect 7300 3337 7308 3343
rect 148 3317 620 3323
rect 628 3317 652 3323
rect 676 3317 700 3323
rect 772 3317 812 3323
rect 1044 3317 1052 3323
rect 1076 3317 1100 3323
rect 1108 3317 1132 3323
rect 1156 3317 1308 3323
rect 1316 3317 1388 3323
rect 1684 3317 1788 3323
rect 1876 3317 2092 3323
rect 2292 3317 2348 3323
rect 2436 3317 2556 3323
rect 3332 3317 3452 3323
rect 3588 3317 3612 3323
rect 3716 3317 3772 3323
rect 3844 3317 3948 3323
rect 4164 3317 4236 3323
rect 4244 3317 4524 3323
rect 4852 3317 5004 3323
rect 5156 3317 5244 3323
rect 5460 3317 5612 3323
rect 6164 3317 6348 3323
rect 6356 3317 6572 3323
rect 6580 3317 6636 3323
rect 6644 3317 6652 3323
rect 6660 3317 6908 3323
rect 6916 3317 7052 3323
rect 7060 3317 7180 3323
rect 7188 3317 7276 3323
rect 7412 3317 7443 3323
rect 116 3297 140 3303
rect 468 3297 508 3303
rect 644 3297 860 3303
rect 1028 3297 1187 3303
rect 1181 3284 1187 3297
rect 1364 3297 1612 3303
rect 1620 3297 1660 3303
rect 1844 3297 1868 3303
rect 1924 3297 1996 3303
rect 2148 3297 2412 3303
rect 2516 3297 2908 3303
rect 3124 3297 3484 3303
rect 3604 3297 3660 3303
rect 3876 3297 3996 3303
rect 4084 3297 4092 3303
rect 4276 3297 4396 3303
rect 4484 3297 4508 3303
rect 4852 3297 5564 3303
rect 5732 3297 6156 3303
rect 6804 3297 6956 3303
rect 7124 3297 7308 3303
rect 180 3277 668 3283
rect 740 3277 940 3283
rect 1012 3277 1084 3283
rect 1092 3277 1148 3283
rect 1188 3277 1324 3283
rect 1588 3277 1836 3283
rect 1972 3277 2012 3283
rect 2036 3277 2060 3283
rect 2212 3277 2636 3283
rect 3092 3277 3404 3283
rect 3412 3277 3548 3283
rect 3556 3277 3724 3283
rect 3892 3277 4060 3283
rect 4340 3277 4572 3283
rect 5124 3277 5164 3283
rect 5172 3277 5244 3283
rect 5252 3277 5532 3283
rect 5572 3277 5660 3283
rect 5668 3277 5676 3283
rect 5780 3277 6476 3283
rect 7204 3277 7276 3283
rect 772 3257 1020 3263
rect 1476 3257 1612 3263
rect 1812 3257 1948 3263
rect 1972 3257 2492 3263
rect 3060 3257 3116 3263
rect 3348 3257 3388 3263
rect 3396 3257 3436 3263
rect 3460 3257 3596 3263
rect 3620 3257 3660 3263
rect 4996 3257 5036 3263
rect 5044 3257 5132 3263
rect 5140 3257 5596 3263
rect 5604 3257 5644 3263
rect 5652 3257 5676 3263
rect 5716 3257 5836 3263
rect 6084 3257 6188 3263
rect 6452 3257 6492 3263
rect 6836 3257 6972 3263
rect 7044 3257 7084 3263
rect 7092 3257 7100 3263
rect 7108 3257 7164 3263
rect 756 3237 876 3243
rect 1284 3237 1580 3243
rect 1748 3237 2444 3243
rect 2468 3237 3100 3243
rect 4628 3237 4876 3243
rect 5460 3237 6044 3243
rect 6596 3237 6668 3243
rect 7213 3243 7219 3256
rect 6996 3237 7219 3243
rect 7284 3237 7356 3243
rect 708 3217 940 3223
rect 1524 3217 1644 3223
rect 1780 3217 2012 3223
rect 2084 3217 2108 3223
rect 2324 3217 2668 3223
rect 3220 3217 3420 3223
rect 5700 3217 5996 3223
rect 7140 3217 7244 3223
rect 1410 3214 1470 3216
rect 1410 3206 1411 3214
rect 1420 3206 1421 3214
rect 1459 3206 1460 3214
rect 1469 3206 1470 3214
rect 1410 3204 1470 3206
rect 4418 3214 4478 3216
rect 4418 3206 4419 3214
rect 4428 3206 4429 3214
rect 4467 3206 4468 3214
rect 4477 3206 4478 3214
rect 4418 3204 4478 3206
rect 772 3197 1372 3203
rect 1540 3197 1708 3203
rect 1732 3197 1836 3203
rect 1940 3197 2140 3203
rect 2356 3197 2732 3203
rect 2788 3197 2828 3203
rect 3316 3197 3628 3203
rect 4036 3197 4140 3203
rect 4740 3197 4780 3203
rect 4788 3197 5436 3203
rect 5652 3197 5772 3203
rect 980 3177 1516 3183
rect 1556 3177 1612 3183
rect 2612 3177 3020 3183
rect 4212 3177 4268 3183
rect 4292 3177 4364 3183
rect 4388 3177 4412 3183
rect 4548 3177 6572 3183
rect 6964 3177 7148 3183
rect 420 3157 812 3163
rect 1156 3157 1244 3163
rect 1524 3157 1564 3163
rect 1940 3157 1948 3163
rect 2388 3157 2444 3163
rect 2548 3157 2828 3163
rect 3012 3157 3052 3163
rect 3460 3157 3740 3163
rect 3780 3157 4588 3163
rect 5396 3157 5612 3163
rect 5620 3157 5820 3163
rect 6468 3157 7260 3163
rect 7268 3157 7340 3163
rect 116 3137 348 3143
rect 804 3137 876 3143
rect 916 3137 1491 3143
rect 212 3117 252 3123
rect 340 3117 396 3123
rect 692 3117 716 3123
rect 724 3117 748 3123
rect 1044 3117 1107 3123
rect 84 3097 204 3103
rect 564 3097 620 3103
rect 820 3097 876 3103
rect 884 3097 908 3103
rect 996 3097 1068 3103
rect 1101 3103 1107 3117
rect 1124 3117 1196 3123
rect 1204 3117 1356 3123
rect 1485 3123 1491 3137
rect 1508 3137 1596 3143
rect 1604 3137 1660 3143
rect 1732 3137 1788 3143
rect 1796 3137 1852 3143
rect 2132 3137 2156 3143
rect 2308 3137 2412 3143
rect 2500 3137 2556 3143
rect 2644 3137 3052 3143
rect 3348 3137 3468 3143
rect 3476 3137 3532 3143
rect 3652 3137 3708 3143
rect 4212 3137 4492 3143
rect 5332 3137 5388 3143
rect 6692 3137 6876 3143
rect 6884 3137 6956 3143
rect 6996 3137 7116 3143
rect 1485 3117 1820 3123
rect 1844 3117 1852 3123
rect 2100 3117 2236 3123
rect 2244 3117 2300 3123
rect 2340 3117 2428 3123
rect 2484 3117 2524 3123
rect 2580 3117 2764 3123
rect 2996 3117 3772 3123
rect 3796 3117 3980 3123
rect 4164 3117 4284 3123
rect 5076 3117 5148 3123
rect 5236 3117 5516 3123
rect 5828 3117 6236 3123
rect 6244 3117 6476 3123
rect 6484 3117 6524 3123
rect 6580 3117 6700 3123
rect 6708 3117 6748 3123
rect 6932 3117 7020 3123
rect 1101 3097 1148 3103
rect 1172 3097 1276 3103
rect 1524 3097 1580 3103
rect 1700 3097 2060 3103
rect 2068 3097 2316 3103
rect 2324 3097 2332 3103
rect 2484 3097 2636 3103
rect 2676 3097 2828 3103
rect 3412 3097 3468 3103
rect 3524 3097 3548 3103
rect 3588 3097 3676 3103
rect 4132 3097 4156 3103
rect 4212 3097 4220 3103
rect 4244 3097 4316 3103
rect 4484 3097 4588 3103
rect 4948 3097 5068 3103
rect 5172 3097 5180 3103
rect 5204 3097 5340 3103
rect 5572 3097 5756 3103
rect 5780 3097 5804 3103
rect 5924 3097 6076 3103
rect 6276 3097 6332 3103
rect 6356 3097 6396 3103
rect 6532 3097 6604 3103
rect 7044 3097 7052 3103
rect 100 3077 268 3083
rect 596 3077 668 3083
rect 724 3077 732 3083
rect 948 3077 1020 3083
rect 1108 3077 1212 3083
rect 1229 3077 1420 3083
rect 84 3057 252 3063
rect 308 3057 364 3063
rect 420 3057 476 3063
rect 516 3057 556 3063
rect 740 3057 764 3063
rect 1229 3063 1235 3077
rect 1428 3077 1884 3083
rect 2020 3077 2380 3083
rect 2548 3077 2588 3083
rect 2676 3077 2796 3083
rect 3412 3077 3628 3083
rect 3652 3077 3980 3083
rect 3997 3083 4003 3096
rect 3997 3077 4140 3083
rect 5204 3077 5372 3083
rect 5508 3077 5724 3083
rect 6180 3077 6188 3083
rect 6292 3077 6300 3083
rect 6468 3077 6556 3083
rect 6564 3077 6636 3083
rect 6644 3077 6860 3083
rect 6884 3077 6956 3083
rect 7316 3077 7340 3083
rect 1044 3057 1235 3063
rect 1284 3057 1500 3063
rect 1540 3057 1932 3063
rect 1940 3057 1964 3063
rect 1972 3057 2108 3063
rect 2116 3057 2220 3063
rect 2228 3057 2284 3063
rect 2548 3057 2588 3063
rect 2980 3057 3036 3063
rect 3444 3057 3596 3063
rect 3732 3057 3788 3063
rect 3828 3057 3852 3063
rect 4100 3057 4204 3063
rect 4308 3057 4332 3063
rect 4340 3057 4348 3063
rect 5172 3057 6076 3063
rect 6084 3057 6204 3063
rect 6324 3057 6588 3063
rect 6820 3057 6924 3063
rect 6996 3057 7084 3063
rect 212 3037 460 3043
rect 644 3037 1148 3043
rect 1524 3037 1644 3043
rect 1652 3037 1708 3043
rect 1716 3037 1772 3043
rect 1780 3037 1804 3043
rect 1812 3037 1836 3043
rect 1876 3037 2508 3043
rect 2532 3037 2780 3043
rect 3300 3037 3500 3043
rect 3716 3037 3788 3043
rect 3988 3037 4204 3043
rect 4244 3037 4364 3043
rect 5060 3037 5164 3043
rect 5444 3037 5484 3043
rect 5492 3037 5580 3043
rect 5588 3037 5628 3043
rect 5860 3037 6092 3043
rect 6132 3037 6364 3043
rect 6372 3037 6460 3043
rect 6484 3037 6652 3043
rect 6660 3037 6908 3043
rect 6916 3037 7052 3043
rect 916 3017 972 3023
rect 1092 3017 1116 3023
rect 1508 3017 1724 3023
rect 1988 3017 2876 3023
rect 3524 3017 3692 3023
rect 3844 3017 4028 3023
rect 4084 3017 4300 3023
rect 4420 3017 4540 3023
rect 4612 3017 4748 3023
rect 5796 3017 5868 3023
rect 6084 3017 6364 3023
rect 6580 3017 6812 3023
rect 6836 3017 7388 3023
rect 2914 3014 2974 3016
rect 2914 3006 2915 3014
rect 2924 3006 2925 3014
rect 2963 3006 2964 3014
rect 2973 3006 2974 3014
rect 2914 3004 2974 3006
rect 5922 3014 5982 3016
rect 5922 3006 5923 3014
rect 5932 3006 5933 3014
rect 5971 3006 5972 3014
rect 5981 3006 5982 3014
rect 5922 3004 5982 3006
rect 820 2997 1196 3003
rect 1364 2997 1580 3003
rect 1828 2997 2380 3003
rect 2404 2997 2428 3003
rect 2708 2997 2748 3003
rect 3220 2997 3644 3003
rect 3716 2997 3772 3003
rect 3908 2997 4172 3003
rect 4212 2997 4300 3003
rect 4372 2997 4604 3003
rect 5108 2997 5260 3003
rect 5460 2997 5900 3003
rect 5997 2997 6300 3003
rect 772 2977 940 2983
rect 948 2977 1196 2983
rect 1652 2977 1868 2983
rect 1908 2977 2140 2983
rect 2196 2977 2396 2983
rect 2564 2977 2812 2983
rect 2884 2977 3132 2983
rect 3428 2977 3484 2983
rect 3492 2977 3724 2983
rect 3732 2977 4012 2983
rect 4020 2977 4156 2983
rect 4164 2977 4412 2983
rect 4820 2977 4876 2983
rect 4884 2977 5196 2983
rect 5220 2977 5292 2983
rect 5997 2983 6003 2997
rect 6340 2997 6540 3003
rect 6708 2997 6844 3003
rect 5316 2977 6003 2983
rect 6196 2977 6620 2983
rect 6788 2977 6972 2983
rect 7012 2977 7052 2983
rect 196 2957 268 2963
rect 500 2957 604 2963
rect 628 2957 716 2963
rect 900 2957 1004 2963
rect 1236 2957 1260 2963
rect 1268 2957 1356 2963
rect 1380 2957 1660 2963
rect 1684 2957 1708 2963
rect 1972 2957 2748 2963
rect 2900 2957 3068 2963
rect 3284 2957 3388 2963
rect 3396 2957 3452 2963
rect 3668 2957 3788 2963
rect 3796 2957 3836 2963
rect 3892 2957 4524 2963
rect 4548 2957 4556 2963
rect 4596 2957 4636 2963
rect 5028 2957 5644 2963
rect 6100 2957 6284 2963
rect 6388 2957 6412 2963
rect 6420 2957 6476 2963
rect 6484 2957 6828 2963
rect 6900 2957 7020 2963
rect 292 2937 364 2943
rect 420 2937 572 2943
rect 580 2937 1020 2943
rect 1156 2937 1212 2943
rect 1220 2937 1468 2943
rect 1572 2937 1676 2943
rect 1748 2937 2012 2943
rect 2020 2937 2028 2943
rect 2036 2937 2108 2943
rect 2244 2937 2300 2943
rect 2900 2937 2940 2943
rect 3236 2937 3356 2943
rect 3476 2937 3612 2943
rect 3620 2937 3676 2943
rect 3700 2937 3740 2943
rect 3748 2937 3932 2943
rect 3940 2937 3996 2943
rect 4004 2937 4188 2943
rect 4196 2937 4316 2943
rect 4340 2937 4508 2943
rect 4900 2937 5052 2943
rect 5236 2937 5340 2943
rect 5412 2937 5500 2943
rect 5828 2937 6252 2943
rect 6628 2937 6988 2943
rect 6996 2937 7068 2943
rect 7076 2937 7244 2943
rect 100 2917 156 2923
rect 212 2917 476 2923
rect 612 2917 636 2923
rect 692 2917 748 2923
rect 820 2917 860 2923
rect 948 2917 1036 2923
rect 1060 2917 1084 2923
rect 1204 2917 1276 2923
rect 1300 2917 1308 2923
rect 1396 2917 1548 2923
rect 1652 2917 1740 2923
rect 1828 2917 1868 2923
rect 1988 2917 2060 2923
rect 2388 2917 2908 2923
rect 3204 2917 3308 2923
rect 3460 2917 3612 2923
rect 3812 2917 3964 2923
rect 4020 2917 4076 2923
rect 4132 2917 4156 2923
rect 4180 2917 4268 2923
rect 4292 2917 4332 2923
rect 4372 2917 4428 2923
rect 4884 2917 4892 2923
rect 5252 2917 5324 2923
rect 5332 2917 5436 2923
rect 5556 2917 5580 2923
rect 5588 2917 6220 2923
rect 6228 2917 6348 2923
rect 6564 2917 6652 2923
rect 7012 2917 7052 2923
rect 7060 2917 7084 2923
rect 7092 2917 7164 2923
rect 596 2897 892 2903
rect 996 2897 1692 2903
rect 1844 2897 2060 2903
rect 2372 2897 2396 2903
rect 2404 2897 2476 2903
rect 2484 2897 2668 2903
rect 2708 2897 2844 2903
rect 3092 2897 3148 2903
rect 3220 2897 3340 2903
rect 3540 2897 3564 2903
rect 3588 2897 3628 2903
rect 3748 2897 3820 2903
rect 3860 2897 3900 2903
rect 3908 2897 4092 2903
rect 4100 2897 4204 2903
rect 4365 2903 4371 2916
rect 4324 2897 4371 2903
rect 4724 2897 5228 2903
rect 5348 2897 5404 2903
rect 5828 2897 5836 2903
rect 5940 2897 5980 2903
rect 5988 2897 6204 2903
rect 6212 2897 6316 2903
rect 6324 2897 6364 2903
rect 6372 2897 6380 2903
rect 6388 2897 6428 2903
rect 6708 2897 6732 2903
rect 6740 2897 7116 2903
rect 388 2877 428 2883
rect 580 2877 668 2883
rect 772 2877 908 2883
rect 1012 2877 1084 2883
rect 1108 2877 1196 2883
rect 1364 2877 1372 2883
rect 1620 2877 1772 2883
rect 2516 2877 2828 2883
rect 2836 2877 2876 2883
rect 3188 2877 3244 2883
rect 3316 2877 3372 2883
rect 3492 2877 3820 2883
rect 3828 2877 3884 2883
rect 3940 2877 4060 2883
rect 4084 2877 4108 2883
rect 4356 2877 4604 2883
rect 5364 2877 5884 2883
rect 5892 2877 6156 2883
rect 6164 2877 6252 2883
rect 6260 2877 6364 2883
rect 6372 2877 6396 2883
rect 6404 2877 6460 2883
rect 6468 2877 6668 2883
rect 6804 2877 6908 2883
rect 244 2857 284 2863
rect 292 2857 364 2863
rect 372 2857 716 2863
rect 1005 2863 1011 2876
rect 724 2857 2044 2863
rect 2052 2857 2204 2863
rect 2212 2857 2284 2863
rect 2292 2857 2300 2863
rect 2308 2857 2444 2863
rect 2452 2857 2540 2863
rect 3268 2857 3356 2863
rect 3933 2863 3939 2876
rect 3364 2857 3939 2863
rect 3956 2857 4252 2863
rect 4276 2857 4412 2863
rect 4628 2857 4748 2863
rect 4756 2857 5020 2863
rect 5236 2857 6140 2863
rect 6516 2857 6604 2863
rect 6612 2857 7187 2863
rect 212 2837 252 2843
rect 260 2837 396 2843
rect 404 2837 668 2843
rect 676 2837 1052 2843
rect 1060 2837 2012 2843
rect 2020 2837 2156 2843
rect 2164 2837 2332 2843
rect 2340 2837 2588 2843
rect 3412 2837 5308 2843
rect 5620 2837 6108 2843
rect 6141 2843 6147 2856
rect 7181 2844 7187 2857
rect 6141 2837 6764 2843
rect 356 2817 492 2823
rect 500 2817 524 2823
rect 532 2817 988 2823
rect 1604 2817 1772 2823
rect 1812 2817 1948 2823
rect 1956 2817 2092 2823
rect 2388 2817 2412 2823
rect 2644 2817 3052 2823
rect 3581 2817 4332 2823
rect 1410 2814 1470 2816
rect 1410 2806 1411 2814
rect 1420 2806 1421 2814
rect 1459 2806 1460 2814
rect 1469 2806 1470 2814
rect 1410 2804 1470 2806
rect 708 2797 780 2803
rect 884 2797 924 2803
rect 932 2797 1100 2803
rect 1252 2797 1292 2803
rect 1540 2797 2771 2803
rect 516 2777 780 2783
rect 884 2777 940 2783
rect 1044 2777 1372 2783
rect 1524 2777 1580 2783
rect 1684 2777 1724 2783
rect 1780 2777 1916 2783
rect 2765 2783 2771 2797
rect 3581 2803 3587 2817
rect 4676 2817 5596 2823
rect 5652 2817 7324 2823
rect 7332 2817 7404 2823
rect 4418 2814 4478 2816
rect 4418 2806 4419 2814
rect 4428 2806 4429 2814
rect 4467 2806 4468 2814
rect 4477 2806 4478 2814
rect 4418 2804 4478 2806
rect 2788 2797 3587 2803
rect 3604 2797 3772 2803
rect 4276 2797 4380 2803
rect 4532 2797 4588 2803
rect 5732 2797 5820 2803
rect 5940 2797 6012 2803
rect 2765 2777 3132 2783
rect 3156 2777 3228 2783
rect 3284 2777 3420 2783
rect 3517 2777 3644 2783
rect 3517 2764 3523 2777
rect 3773 2783 3779 2796
rect 3773 2777 3980 2783
rect 4420 2777 4844 2783
rect 5332 2777 5388 2783
rect 6308 2777 6332 2783
rect 6340 2777 6924 2783
rect 468 2757 652 2763
rect 804 2757 860 2763
rect 1028 2757 1340 2763
rect 1348 2757 1644 2763
rect 1668 2757 1868 2763
rect 1908 2757 1948 2763
rect 2676 2757 2700 2763
rect 3380 2757 3516 2763
rect 3556 2757 3596 2763
rect 3684 2757 3724 2763
rect 3748 2757 3868 2763
rect 3972 2757 4044 2763
rect 4180 2757 4652 2763
rect 5444 2757 5788 2763
rect 5812 2757 6028 2763
rect 7348 2757 7404 2763
rect 404 2737 444 2743
rect 596 2737 620 2743
rect 660 2737 748 2743
rect 756 2737 1500 2743
rect 1508 2737 1708 2743
rect 1716 2737 2252 2743
rect 2868 2737 3571 2743
rect 516 2717 764 2723
rect 820 2717 892 2723
rect 900 2717 1804 2723
rect 1812 2717 2140 2723
rect 2148 2717 2220 2723
rect 2228 2717 2396 2723
rect 2404 2717 2444 2723
rect 2564 2717 2652 2723
rect 3252 2717 3420 2723
rect 3508 2717 3548 2723
rect 3565 2723 3571 2737
rect 3588 2737 3788 2743
rect 3796 2737 3804 2743
rect 3844 2737 4060 2743
rect 4084 2737 4092 2743
rect 4116 2737 4236 2743
rect 4308 2737 4492 2743
rect 4500 2737 4556 2743
rect 5108 2737 5484 2743
rect 5588 2737 5772 2743
rect 5780 2737 5900 2743
rect 5908 2737 6108 2743
rect 6404 2737 6716 2743
rect 6772 2737 6892 2743
rect 6932 2737 7004 2743
rect 3565 2717 3676 2723
rect 3732 2717 4156 2723
rect 4196 2717 4364 2723
rect 4372 2717 4604 2723
rect 5076 2717 5148 2723
rect 5236 2717 5708 2723
rect 5716 2717 5772 2723
rect 5796 2717 6204 2723
rect 6612 2717 6796 2723
rect 6980 2717 7068 2723
rect 7092 2717 7148 2723
rect 7156 2717 7340 2723
rect 100 2697 300 2703
rect 564 2697 1004 2703
rect 1012 2697 1132 2703
rect 1156 2697 1164 2703
rect 1172 2697 1180 2703
rect 1268 2697 1388 2703
rect 1572 2697 1580 2703
rect 1652 2697 1676 2703
rect 1716 2697 1756 2703
rect 2116 2697 2268 2703
rect 2692 2697 2716 2703
rect 2788 2697 2860 2703
rect 3204 2697 3260 2703
rect 3364 2697 3596 2703
rect 3732 2697 4019 2703
rect 340 2677 364 2683
rect 548 2677 956 2683
rect 1028 2677 1068 2683
rect 1076 2677 1164 2683
rect 1204 2677 1276 2683
rect 1284 2677 1868 2683
rect 1876 2677 2412 2683
rect 2548 2677 2572 2683
rect 2660 2677 2716 2683
rect 2772 2677 2876 2683
rect 3108 2677 3212 2683
rect 3332 2677 3356 2683
rect 3428 2677 3916 2683
rect 3924 2677 3996 2683
rect 4013 2683 4019 2697
rect 4148 2697 4156 2703
rect 4180 2697 4204 2703
rect 4221 2697 4803 2703
rect 4221 2683 4227 2697
rect 4013 2677 4227 2683
rect 4276 2677 4611 2683
rect 244 2657 332 2663
rect 724 2657 828 2663
rect 916 2657 1004 2663
rect 1236 2657 1324 2663
rect 1332 2657 1660 2663
rect 1684 2657 1955 2663
rect 324 2637 572 2643
rect 868 2637 972 2643
rect 1092 2637 1148 2643
rect 1188 2637 1244 2643
rect 1252 2637 1299 2643
rect 372 2617 1244 2623
rect 1293 2623 1299 2637
rect 1316 2637 1852 2643
rect 1860 2637 1900 2643
rect 1949 2643 1955 2657
rect 1972 2657 1996 2663
rect 2404 2657 2476 2663
rect 2740 2657 2828 2663
rect 3220 2657 3276 2663
rect 3540 2657 3564 2663
rect 3668 2657 3708 2663
rect 3844 2657 3852 2663
rect 4020 2657 4108 2663
rect 4164 2657 4204 2663
rect 4260 2657 4300 2663
rect 4308 2657 4540 2663
rect 4564 2657 4588 2663
rect 4605 2663 4611 2677
rect 4644 2677 4780 2683
rect 4797 2683 4803 2697
rect 4852 2697 4876 2703
rect 4884 2697 5004 2703
rect 5156 2697 5164 2703
rect 5172 2697 5196 2703
rect 5204 2697 5340 2703
rect 5508 2697 5548 2703
rect 5716 2697 5756 2703
rect 6004 2697 6140 2703
rect 6276 2697 6460 2703
rect 6612 2697 6876 2703
rect 6884 2697 6972 2703
rect 7348 2697 7356 2703
rect 4797 2677 4956 2683
rect 5412 2677 5468 2683
rect 5556 2677 5644 2683
rect 5748 2677 5868 2683
rect 5876 2677 6028 2683
rect 6132 2677 6172 2683
rect 6196 2677 6284 2683
rect 6292 2677 6316 2683
rect 6436 2677 6460 2683
rect 6532 2677 6892 2683
rect 7172 2677 7196 2683
rect 7204 2677 7244 2683
rect 4605 2657 5212 2663
rect 5380 2657 5436 2663
rect 5492 2657 5804 2663
rect 5828 2657 5868 2663
rect 5885 2657 6396 2663
rect 1949 2637 2060 2643
rect 2228 2637 2284 2643
rect 2468 2637 2540 2643
rect 3204 2637 3404 2643
rect 3684 2637 3900 2643
rect 4004 2637 4924 2643
rect 4964 2637 5820 2643
rect 5885 2643 5891 2657
rect 6500 2657 6556 2663
rect 6564 2657 6684 2663
rect 6852 2657 7116 2663
rect 5860 2637 5891 2643
rect 6260 2637 6316 2643
rect 6372 2637 6636 2643
rect 6756 2637 7020 2643
rect 1293 2617 1788 2623
rect 2052 2617 2204 2623
rect 2340 2617 2396 2623
rect 3092 2617 3196 2623
rect 3444 2617 4268 2623
rect 4292 2617 4636 2623
rect 4724 2617 4828 2623
rect 4948 2617 5020 2623
rect 5028 2617 5196 2623
rect 5380 2617 5788 2623
rect 5828 2617 5836 2623
rect 6068 2617 6140 2623
rect 6420 2617 6508 2623
rect 6516 2617 6876 2623
rect 6884 2617 6924 2623
rect 7060 2617 7132 2623
rect 2914 2614 2974 2616
rect 2914 2606 2915 2614
rect 2924 2606 2925 2614
rect 2963 2606 2964 2614
rect 2973 2606 2974 2614
rect 2914 2604 2974 2606
rect 5922 2614 5982 2616
rect 5922 2606 5923 2614
rect 5932 2606 5933 2614
rect 5971 2606 5972 2614
rect 5981 2606 5982 2614
rect 5922 2604 5982 2606
rect 964 2597 2124 2603
rect 2132 2597 2156 2603
rect 2164 2597 2364 2603
rect 2372 2597 2508 2603
rect 3124 2597 3148 2603
rect 3652 2597 3884 2603
rect 3924 2597 3948 2603
rect 3988 2597 4076 2603
rect 4100 2597 4108 2603
rect 4132 2597 4140 2603
rect 4228 2597 4252 2603
rect 4580 2597 4876 2603
rect 5236 2597 5516 2603
rect 5748 2597 5804 2603
rect 6132 2597 6620 2603
rect 6772 2597 6860 2603
rect 6868 2597 6988 2603
rect 7012 2597 7036 2603
rect 836 2577 1548 2583
rect 1556 2577 1612 2583
rect 1844 2577 2204 2583
rect 2500 2577 3020 2583
rect 3124 2577 3148 2583
rect 3332 2577 3772 2583
rect 3796 2577 3868 2583
rect 3988 2577 4076 2583
rect 4132 2577 4284 2583
rect 4516 2577 4620 2583
rect 4692 2577 4716 2583
rect 4740 2577 4764 2583
rect 4788 2577 4940 2583
rect 5284 2577 6444 2583
rect 6548 2577 6588 2583
rect 6740 2577 6748 2583
rect 6884 2577 6988 2583
rect 7108 2577 7148 2583
rect 7188 2577 7372 2583
rect 404 2557 460 2563
rect 676 2557 700 2563
rect 1092 2557 1164 2563
rect 1300 2557 1324 2563
rect 1428 2557 1548 2563
rect 1556 2557 1628 2563
rect 1732 2557 1756 2563
rect 1821 2563 1827 2576
rect 1821 2557 1868 2563
rect 1940 2557 1980 2563
rect 2036 2557 2092 2563
rect 2292 2557 2428 2563
rect 3284 2557 3564 2563
rect 3588 2557 3644 2563
rect 3668 2557 3740 2563
rect 3764 2557 3788 2563
rect 3812 2557 3836 2563
rect 3876 2557 3916 2563
rect 3940 2557 3980 2563
rect 3988 2557 4028 2563
rect 4068 2557 4092 2563
rect 4116 2557 4540 2563
rect 4596 2557 4700 2563
rect 4708 2557 4812 2563
rect 4820 2557 5004 2563
rect 5460 2557 5516 2563
rect 5540 2557 5692 2563
rect 5812 2557 6124 2563
rect 6308 2557 6684 2563
rect 212 2537 236 2543
rect 324 2537 380 2543
rect 388 2537 460 2543
rect 468 2537 508 2543
rect 1284 2537 1308 2543
rect 1572 2537 1596 2543
rect 1748 2537 1852 2543
rect 1908 2537 1948 2543
rect 2020 2537 2380 2543
rect 2836 2537 2860 2543
rect 3380 2537 3628 2543
rect 3636 2537 3660 2543
rect 3684 2537 3820 2543
rect 3828 2537 3916 2543
rect 3924 2537 4188 2543
rect 4244 2537 4371 2543
rect 68 2517 204 2523
rect 212 2517 540 2523
rect 596 2517 636 2523
rect 772 2517 828 2523
rect 932 2517 1052 2523
rect 1140 2517 1180 2523
rect 1348 2517 1388 2523
rect 1860 2517 1884 2523
rect 2004 2517 2236 2523
rect 2708 2517 2716 2523
rect 2804 2517 2844 2523
rect 3076 2517 3100 2523
rect 3508 2517 3564 2523
rect 3732 2517 3820 2523
rect 3828 2517 3868 2523
rect 3972 2517 4028 2523
rect 4052 2517 4172 2523
rect 4205 2517 4332 2523
rect 116 2497 252 2503
rect 260 2497 588 2503
rect 596 2497 892 2503
rect 1204 2497 1308 2503
rect 1332 2497 1436 2503
rect 1524 2497 1548 2503
rect 1636 2497 2188 2503
rect 2196 2497 2204 2503
rect 2228 2497 2332 2503
rect 2452 2497 2476 2503
rect 2820 2497 2844 2503
rect 3300 2497 3436 2503
rect 3636 2497 3676 2503
rect 3764 2497 4076 2503
rect 4084 2497 4092 2503
rect 4205 2503 4211 2517
rect 4365 2523 4371 2537
rect 4532 2537 4652 2543
rect 4692 2537 4700 2543
rect 4740 2537 4780 2543
rect 5556 2537 5852 2543
rect 5860 2537 6028 2543
rect 6036 2537 6108 2543
rect 6372 2537 6492 2543
rect 6516 2537 6556 2543
rect 4365 2517 4508 2523
rect 4564 2517 4572 2523
rect 4692 2517 4732 2523
rect 4772 2517 4908 2523
rect 5316 2517 5580 2523
rect 5652 2517 5900 2523
rect 6020 2517 6028 2523
rect 6036 2517 6364 2523
rect 6388 2517 6444 2523
rect 6740 2517 6812 2523
rect 6868 2517 6956 2523
rect 6909 2504 6915 2517
rect 7284 2517 7292 2523
rect 4116 2497 4211 2503
rect 4228 2497 4268 2503
rect 4468 2497 4508 2503
rect 4596 2497 4604 2503
rect 4852 2497 4860 2503
rect 5412 2497 5564 2503
rect 5572 2497 5612 2503
rect 5988 2497 6428 2503
rect 6452 2497 6492 2503
rect 6660 2497 6812 2503
rect 6852 2497 6908 2503
rect 6964 2497 7100 2503
rect 340 2477 396 2483
rect 404 2477 444 2483
rect 452 2477 524 2483
rect 532 2477 684 2483
rect 788 2477 1884 2483
rect 1924 2477 2028 2483
rect 2132 2477 2156 2483
rect 2244 2477 2764 2483
rect 3700 2477 4012 2483
rect 4020 2477 4252 2483
rect 4308 2477 4524 2483
rect 4644 2477 5340 2483
rect 5396 2477 5644 2483
rect 5652 2477 5740 2483
rect 5780 2477 6028 2483
rect 6100 2477 6252 2483
rect 6964 2477 6972 2483
rect 1236 2457 1420 2463
rect 1444 2457 1580 2463
rect 1588 2457 1996 2463
rect 2020 2457 2204 2463
rect 2212 2457 2268 2463
rect 2397 2457 2787 2463
rect 612 2437 1532 2443
rect 1588 2437 1612 2443
rect 2397 2443 2403 2457
rect 1748 2437 2403 2443
rect 2420 2437 2700 2443
rect 2781 2443 2787 2457
rect 2804 2457 4108 2463
rect 4148 2457 4291 2463
rect 4285 2444 4291 2457
rect 4372 2457 4412 2463
rect 4532 2457 4716 2463
rect 4868 2457 5132 2463
rect 5140 2457 5404 2463
rect 5428 2457 5500 2463
rect 5508 2457 5596 2463
rect 5604 2457 5772 2463
rect 5812 2457 6140 2463
rect 6452 2457 6876 2463
rect 2781 2437 2972 2443
rect 3364 2437 3484 2443
rect 3492 2437 3516 2443
rect 3604 2437 3756 2443
rect 3780 2437 3868 2443
rect 3885 2437 4252 2443
rect 1012 2417 1100 2423
rect 1188 2417 1324 2423
rect 1748 2417 1772 2423
rect 1908 2417 2604 2423
rect 3396 2417 3452 2423
rect 3476 2417 3724 2423
rect 3885 2423 3891 2437
rect 4292 2437 4780 2443
rect 5492 2437 5868 2443
rect 5876 2437 6540 2443
rect 6708 2437 7260 2443
rect 3780 2417 3891 2423
rect 3908 2417 4044 2423
rect 4100 2417 4204 2423
rect 4228 2417 4300 2423
rect 4676 2417 4908 2423
rect 5332 2417 5484 2423
rect 5492 2417 5580 2423
rect 5780 2417 5836 2423
rect 6484 2417 6700 2423
rect 1410 2414 1470 2416
rect 1410 2406 1411 2414
rect 1420 2406 1421 2414
rect 1459 2406 1460 2414
rect 1469 2406 1470 2414
rect 1410 2404 1470 2406
rect 4418 2414 4478 2416
rect 4418 2406 4419 2414
rect 4428 2406 4429 2414
rect 4467 2406 4468 2414
rect 4477 2406 4478 2414
rect 4418 2404 4478 2406
rect 1252 2397 1395 2403
rect 532 2377 1004 2383
rect 1092 2377 1196 2383
rect 1204 2377 1212 2383
rect 1220 2377 1244 2383
rect 1389 2383 1395 2397
rect 1892 2397 2988 2403
rect 3204 2397 3692 2403
rect 3828 2397 3916 2403
rect 4020 2397 4236 2403
rect 4260 2397 4396 2403
rect 4548 2397 4716 2403
rect 5204 2397 5404 2403
rect 6468 2397 6620 2403
rect 6708 2397 7180 2403
rect 1389 2377 1740 2383
rect 1764 2377 2572 2383
rect 2580 2377 2780 2383
rect 3028 2377 4188 2383
rect 4212 2377 4700 2383
rect 5284 2377 5372 2383
rect 5428 2377 5612 2383
rect 5892 2377 6044 2383
rect 6068 2377 6076 2383
rect 6084 2377 6316 2383
rect 6420 2377 6700 2383
rect 6868 2377 7212 2383
rect 180 2357 492 2363
rect 500 2357 668 2363
rect 1044 2357 1244 2363
rect 1524 2357 1932 2363
rect 2500 2357 2748 2363
rect 3012 2357 3052 2363
rect 3588 2357 3708 2363
rect 3716 2357 3884 2363
rect 4052 2357 4076 2363
rect 4132 2357 4252 2363
rect 4500 2357 4540 2363
rect 4564 2357 4620 2363
rect 4644 2357 5100 2363
rect 5156 2357 5484 2363
rect 5716 2357 6956 2363
rect 6964 2357 7372 2363
rect 388 2337 428 2343
rect 580 2337 620 2343
rect 772 2337 780 2343
rect 916 2337 972 2343
rect 1124 2337 1532 2343
rect 1556 2337 1692 2343
rect 1700 2337 1788 2343
rect 1796 2337 1804 2343
rect 2164 2337 2268 2343
rect 2308 2337 2508 2343
rect 2788 2337 3084 2343
rect 3124 2337 3148 2343
rect 3284 2337 3596 2343
rect 3645 2337 3740 2343
rect 3645 2324 3651 2337
rect 3748 2337 3900 2343
rect 3917 2337 3964 2343
rect 116 2317 236 2323
rect 468 2317 540 2323
rect 660 2317 1020 2323
rect 1172 2317 1228 2323
rect 1428 2317 1580 2323
rect 1668 2317 1964 2323
rect 2052 2317 2124 2323
rect 2260 2317 2268 2323
rect 2548 2317 2668 2323
rect 2676 2317 3116 2323
rect 3172 2317 3244 2323
rect 3380 2317 3612 2323
rect 3661 2317 3772 2323
rect 148 2297 284 2303
rect 340 2297 364 2303
rect 461 2297 620 2303
rect 461 2284 467 2297
rect 692 2297 716 2303
rect 772 2297 828 2303
rect 836 2297 876 2303
rect 916 2297 1132 2303
rect 1140 2297 1260 2303
rect 1284 2297 1308 2303
rect 1348 2297 1356 2303
rect 1476 2297 1900 2303
rect 1908 2297 2092 2303
rect 2276 2297 2316 2303
rect 2756 2297 2780 2303
rect 2788 2297 2860 2303
rect 2868 2297 3020 2303
rect 3028 2297 3084 2303
rect 3092 2297 3148 2303
rect 3156 2297 3276 2303
rect 3508 2297 3523 2303
rect 100 2277 428 2283
rect 436 2277 460 2283
rect 532 2277 572 2283
rect 740 2277 764 2283
rect 788 2277 844 2283
rect 852 2277 972 2283
rect 980 2277 1052 2283
rect 1300 2277 1340 2283
rect 1460 2277 1660 2283
rect 1668 2277 1724 2283
rect 1732 2277 1772 2283
rect 1844 2277 1868 2283
rect 1908 2277 2044 2283
rect 2116 2277 2140 2283
rect 2356 2277 2396 2283
rect 2516 2277 2556 2283
rect 2756 2277 2764 2283
rect 2772 2277 2796 2283
rect 2820 2277 3020 2283
rect 3044 2277 3100 2283
rect 3108 2277 3164 2283
rect 3172 2277 3292 2283
rect 3517 2283 3523 2297
rect 3540 2297 3548 2303
rect 3556 2297 3564 2303
rect 3661 2303 3667 2317
rect 3917 2323 3923 2337
rect 4084 2337 4492 2343
rect 4500 2337 5052 2343
rect 5204 2337 5692 2343
rect 5700 2337 5804 2343
rect 5844 2337 6540 2343
rect 6772 2337 6972 2343
rect 3876 2317 3923 2323
rect 3940 2317 3996 2323
rect 4020 2317 4428 2323
rect 4436 2317 4588 2323
rect 4596 2317 4652 2323
rect 4660 2317 4716 2323
rect 4820 2317 5308 2323
rect 5380 2317 5468 2323
rect 5508 2317 5612 2323
rect 5668 2317 5788 2323
rect 5812 2317 6108 2323
rect 6116 2317 6156 2323
rect 6308 2317 6380 2323
rect 6500 2317 6556 2323
rect 6564 2317 6572 2323
rect 6868 2317 6940 2323
rect 3604 2297 3667 2303
rect 3684 2297 3756 2303
rect 3821 2297 3980 2303
rect 3517 2277 3548 2283
rect 3636 2277 3692 2283
rect 3821 2283 3827 2297
rect 4052 2297 4268 2303
rect 4276 2297 4316 2303
rect 4404 2297 4691 2303
rect 3716 2277 3827 2283
rect 3844 2277 3884 2283
rect 3892 2277 3948 2283
rect 3972 2277 4108 2283
rect 4180 2277 4556 2283
rect 4564 2277 4588 2283
rect 4644 2277 4652 2283
rect 4685 2283 4691 2297
rect 4708 2297 4716 2303
rect 4756 2297 5052 2303
rect 5124 2297 5212 2303
rect 5236 2297 5324 2303
rect 5348 2297 5388 2303
rect 5396 2297 5564 2303
rect 5620 2297 5788 2303
rect 5812 2297 5939 2303
rect 4685 2277 4844 2283
rect 5060 2277 5084 2283
rect 5188 2277 5292 2283
rect 5364 2277 5500 2283
rect 5652 2277 5676 2283
rect 5716 2277 5740 2283
rect 5764 2277 5916 2283
rect 5933 2283 5939 2297
rect 6100 2297 6156 2303
rect 6164 2297 6220 2303
rect 6244 2297 6284 2303
rect 6340 2297 6444 2303
rect 6468 2297 6572 2303
rect 6580 2297 6636 2303
rect 6660 2297 6684 2303
rect 6820 2297 6892 2303
rect 6900 2297 6940 2303
rect 7316 2297 7372 2303
rect 5933 2277 6188 2283
rect 6205 2277 6380 2283
rect 20 2257 124 2263
rect 468 2257 492 2263
rect 884 2257 1164 2263
rect 1172 2257 1212 2263
rect 1300 2257 1340 2263
rect 1517 2257 1740 2263
rect 868 2237 908 2243
rect 1028 2237 1100 2243
rect 1517 2243 1523 2257
rect 1748 2257 1852 2263
rect 2388 2257 2428 2263
rect 2548 2257 2572 2263
rect 2612 2257 2668 2263
rect 2676 2257 2684 2263
rect 3476 2257 3532 2263
rect 3668 2257 3852 2263
rect 3956 2257 3996 2263
rect 4164 2257 4204 2263
rect 4221 2257 4732 2263
rect 1316 2237 1523 2243
rect 1540 2237 2492 2243
rect 2852 2237 2860 2243
rect 2916 2237 3228 2243
rect 3268 2237 3308 2243
rect 3348 2237 3372 2243
rect 3380 2237 3596 2243
rect 3636 2237 3660 2243
rect 3700 2237 3740 2243
rect 3780 2237 3868 2243
rect 3924 2237 4060 2243
rect 4221 2243 4227 2257
rect 4804 2257 5491 2263
rect 4196 2237 4227 2243
rect 4237 2237 4300 2243
rect 852 2217 956 2223
rect 1140 2217 1468 2223
rect 2532 2217 2604 2223
rect 2628 2217 2732 2223
rect 3236 2217 3532 2223
rect 3540 2217 3660 2223
rect 3757 2223 3763 2236
rect 4237 2224 4243 2237
rect 4324 2237 4355 2243
rect 3757 2217 3948 2223
rect 4036 2217 4156 2223
rect 4164 2217 4236 2223
rect 4308 2217 4332 2223
rect 4349 2223 4355 2237
rect 4580 2237 4684 2243
rect 5076 2237 5148 2243
rect 5444 2237 5468 2243
rect 5485 2243 5491 2257
rect 5508 2257 5532 2263
rect 5588 2257 5692 2263
rect 5732 2257 5772 2263
rect 5828 2257 6060 2263
rect 6205 2263 6211 2277
rect 6564 2277 6668 2283
rect 6900 2277 7116 2283
rect 6180 2257 6211 2263
rect 6372 2257 6652 2263
rect 6804 2257 6924 2263
rect 5485 2237 6508 2243
rect 6532 2237 6604 2243
rect 6724 2237 6844 2243
rect 6980 2237 7404 2243
rect 4349 2217 4748 2223
rect 4964 2217 5116 2223
rect 5380 2217 5708 2223
rect 5748 2217 5868 2223
rect 6068 2217 6220 2223
rect 6244 2217 6588 2223
rect 6596 2217 6851 2223
rect 2914 2214 2974 2216
rect 2914 2206 2915 2214
rect 2924 2206 2925 2214
rect 2963 2206 2964 2214
rect 2973 2206 2974 2214
rect 2914 2204 2974 2206
rect 5922 2214 5982 2216
rect 5922 2206 5923 2214
rect 5932 2206 5933 2214
rect 5971 2206 5972 2214
rect 5981 2206 5982 2214
rect 5922 2204 5982 2206
rect 6845 2204 6851 2217
rect 7108 2217 7132 2223
rect 7172 2217 7180 2223
rect 1204 2197 2796 2203
rect 3412 2197 3436 2203
rect 3460 2197 3692 2203
rect 3940 2197 4012 2203
rect 4116 2197 4620 2203
rect 4836 2197 5180 2203
rect 5684 2197 5836 2203
rect 6148 2197 6172 2203
rect 6628 2197 6668 2203
rect 6692 2197 6732 2203
rect 6852 2197 6924 2203
rect 6996 2197 7052 2203
rect 500 2177 988 2183
rect 1076 2177 1628 2183
rect 1796 2177 1852 2183
rect 1860 2177 1900 2183
rect 1924 2177 2076 2183
rect 2116 2177 2140 2183
rect 2196 2177 2620 2183
rect 2644 2177 2684 2183
rect 2756 2177 3036 2183
rect 3412 2177 3612 2183
rect 3780 2177 3836 2183
rect 3844 2177 3980 2183
rect 4004 2177 4268 2183
rect 4292 2177 4524 2183
rect 4541 2177 4668 2183
rect 276 2157 652 2163
rect 1284 2157 1340 2163
rect 1364 2157 1404 2163
rect 1780 2157 2028 2163
rect 2100 2157 2316 2163
rect 2468 2157 2540 2163
rect 2676 2157 2748 2163
rect 3124 2157 3452 2163
rect 3476 2157 3516 2163
rect 3572 2157 4076 2163
rect 4100 2157 4124 2163
rect 4148 2157 4188 2163
rect 4260 2157 4364 2163
rect 4541 2163 4547 2177
rect 4676 2177 4940 2183
rect 4980 2177 5628 2183
rect 5652 2177 5756 2183
rect 5972 2177 6268 2183
rect 6276 2177 6316 2183
rect 6372 2177 6412 2183
rect 6420 2177 6556 2183
rect 6932 2177 6940 2183
rect 7204 2177 7340 2183
rect 4516 2157 4547 2163
rect 4589 2157 5004 2163
rect 4589 2144 4595 2157
rect 5588 2157 5660 2163
rect 5668 2157 5772 2163
rect 6036 2157 6204 2163
rect 6228 2157 6636 2163
rect 6900 2157 6988 2163
rect 212 2137 316 2143
rect 452 2137 684 2143
rect 756 2137 828 2143
rect 900 2137 940 2143
rect 948 2137 1004 2143
rect 1012 2137 1068 2143
rect 1076 2137 1132 2143
rect 1332 2137 1964 2143
rect 2052 2137 2252 2143
rect 2340 2137 2460 2143
rect 2468 2137 2572 2143
rect 2788 2137 2956 2143
rect 3124 2137 3228 2143
rect 3316 2137 3372 2143
rect 3380 2137 3468 2143
rect 3476 2137 3484 2143
rect 3492 2137 3500 2143
rect 3508 2137 3580 2143
rect 3604 2137 3852 2143
rect 3860 2137 4364 2143
rect 4548 2137 4588 2143
rect 4612 2137 4716 2143
rect 4884 2137 5004 2143
rect 5332 2137 5404 2143
rect 5620 2137 5868 2143
rect 5940 2137 6124 2143
rect 6260 2137 6348 2143
rect 6356 2137 6588 2143
rect 6788 2137 6908 2143
rect 6916 2137 6956 2143
rect 7092 2137 7116 2143
rect 52 2117 252 2123
rect 308 2117 380 2123
rect 436 2117 476 2123
rect 516 2117 524 2123
rect 548 2117 652 2123
rect 804 2117 1308 2123
rect 1364 2117 1516 2123
rect 1700 2117 2115 2123
rect 180 2097 284 2103
rect 404 2097 620 2103
rect 628 2097 924 2103
rect 932 2097 1228 2103
rect 1236 2097 1244 2103
rect 1412 2097 1516 2103
rect 1604 2097 1676 2103
rect 1700 2097 1852 2103
rect 1940 2097 1964 2103
rect 2109 2103 2115 2117
rect 2212 2117 2268 2123
rect 2308 2117 2364 2123
rect 2372 2117 2668 2123
rect 2724 2117 2828 2123
rect 3028 2117 3164 2123
rect 3172 2117 3212 2123
rect 3252 2117 3260 2123
rect 3636 2117 3644 2123
rect 3732 2117 3772 2123
rect 4020 2117 4028 2123
rect 4148 2117 4236 2123
rect 4260 2117 4268 2123
rect 4356 2117 4492 2123
rect 4644 2117 4652 2123
rect 5012 2117 5052 2123
rect 5060 2117 5164 2123
rect 5188 2117 5260 2123
rect 5268 2117 5356 2123
rect 5492 2117 5580 2123
rect 5652 2117 5676 2123
rect 5924 2117 5980 2123
rect 6100 2117 6140 2123
rect 6276 2117 6444 2123
rect 6468 2117 6508 2123
rect 6516 2117 6620 2123
rect 6628 2117 6828 2123
rect 6836 2117 6860 2123
rect 6884 2117 7036 2123
rect 7060 2117 7084 2123
rect 7124 2117 7148 2123
rect 2109 2097 2188 2103
rect 2260 2097 2428 2103
rect 2548 2097 2556 2103
rect 2804 2097 2867 2103
rect 2861 2084 2867 2097
rect 3124 2097 3836 2103
rect 3876 2097 3932 2103
rect 4020 2097 4044 2103
rect 4052 2097 4204 2103
rect 4308 2097 4348 2103
rect 4372 2097 4396 2103
rect 4484 2097 4604 2103
rect 4772 2097 4796 2103
rect 5524 2097 5564 2103
rect 5572 2097 5884 2103
rect 6180 2097 6572 2103
rect 6724 2097 6764 2103
rect 6772 2097 7116 2103
rect 7124 2097 7292 2103
rect 100 2077 172 2083
rect 212 2077 316 2083
rect 324 2077 540 2083
rect 676 2077 700 2083
rect 820 2077 876 2083
rect 932 2077 988 2083
rect 996 2077 1052 2083
rect 1060 2077 1116 2083
rect 1213 2077 1564 2083
rect 148 2057 172 2063
rect 532 2057 556 2063
rect 740 2057 940 2063
rect 1213 2063 1219 2077
rect 1572 2077 1628 2083
rect 1684 2077 1708 2083
rect 1716 2077 1772 2083
rect 1812 2077 2844 2083
rect 3076 2077 4012 2083
rect 4036 2077 4060 2083
rect 4084 2077 4316 2083
rect 4420 2077 4684 2083
rect 5252 2077 5260 2083
rect 5268 2077 5292 2083
rect 5300 2077 5772 2083
rect 5908 2077 6060 2083
rect 6164 2077 6172 2083
rect 6340 2077 6684 2083
rect 7060 2077 7164 2083
rect 980 2057 1219 2063
rect 1316 2057 1436 2063
rect 1572 2057 1612 2063
rect 1860 2057 1916 2063
rect 2004 2057 2060 2063
rect 2180 2057 2236 2063
rect 2324 2057 2364 2063
rect 2388 2057 2412 2063
rect 2452 2057 2508 2063
rect 3460 2057 4780 2063
rect 5108 2057 5148 2063
rect 5156 2057 5596 2063
rect 5796 2057 6780 2063
rect 356 2037 588 2043
rect 724 2037 732 2043
rect 1236 2037 1324 2043
rect 1389 2037 1708 2043
rect 1389 2023 1395 2037
rect 1796 2037 2028 2043
rect 2084 2037 2380 2043
rect 2404 2037 3212 2043
rect 3380 2037 3548 2043
rect 3556 2037 3596 2043
rect 3684 2037 3724 2043
rect 3764 2037 3804 2043
rect 4036 2037 4508 2043
rect 4708 2037 4876 2043
rect 4916 2037 5068 2043
rect 5332 2037 5484 2043
rect 6100 2037 6124 2043
rect 6164 2037 6540 2043
rect 6820 2037 6828 2043
rect 7172 2037 7180 2043
rect 1140 2017 1395 2023
rect 1604 2017 1644 2023
rect 1876 2017 1916 2023
rect 2196 2017 2460 2023
rect 2516 2017 2668 2023
rect 2852 2017 3372 2023
rect 3396 2017 3580 2023
rect 3796 2017 4220 2023
rect 4244 2017 4380 2023
rect 4980 2017 5100 2023
rect 5348 2017 5660 2023
rect 5668 2017 6076 2023
rect 6292 2017 6300 2023
rect 6340 2017 7180 2023
rect 7188 2017 7340 2023
rect 1410 2014 1470 2016
rect 1410 2006 1411 2014
rect 1420 2006 1421 2014
rect 1459 2006 1460 2014
rect 1469 2006 1470 2014
rect 1410 2004 1470 2006
rect 4418 2014 4478 2016
rect 4418 2006 4419 2014
rect 4428 2006 4429 2014
rect 4467 2006 4468 2014
rect 4477 2006 4478 2014
rect 4418 2004 4478 2006
rect 356 1997 1196 2003
rect 1300 1997 1372 2003
rect 2116 1997 2316 2003
rect 2340 1997 2876 2003
rect 2884 1997 3052 2003
rect 3060 1997 3276 2003
rect 3284 1997 3436 2003
rect 3444 1997 3756 2003
rect 3764 1997 3788 2003
rect 3972 1997 4060 2003
rect 4132 1997 4252 2003
rect 4996 1997 5052 2003
rect 5060 1997 5420 2003
rect 5428 1997 5740 2003
rect 6052 1997 6108 2003
rect 6116 1997 6236 2003
rect 6244 1997 6428 2003
rect 6548 1997 7116 2003
rect 7188 1997 7228 2003
rect 708 1977 780 1983
rect 1332 1977 1356 1983
rect 1380 1977 1548 1983
rect 1556 1977 1836 1983
rect 1844 1977 1900 1983
rect 1924 1977 2764 1983
rect 3236 1977 3340 1983
rect 3364 1977 4380 1983
rect 4404 1977 4444 1983
rect 4468 1977 4572 1983
rect 5076 1977 5340 1983
rect 5348 1977 5372 1983
rect 5396 1977 5580 1983
rect 5796 1977 6028 1983
rect 6100 1977 6620 1983
rect 6676 1977 6844 1983
rect 1284 1957 1308 1963
rect 1348 1957 1388 1963
rect 1396 1957 1564 1963
rect 1572 1957 1580 1963
rect 1588 1957 1612 1963
rect 1620 1957 1676 1963
rect 1684 1957 1724 1963
rect 1732 1957 1852 1963
rect 1860 1957 1916 1963
rect 2356 1957 2780 1963
rect 2820 1957 3276 1963
rect 3348 1957 3564 1963
rect 3732 1957 4172 1963
rect 4196 1957 4284 1963
rect 4340 1957 4540 1963
rect 4548 1957 4604 1963
rect 4612 1957 4828 1963
rect 5556 1957 5708 1963
rect 5716 1957 5932 1963
rect 5940 1957 6156 1963
rect 6164 1957 6412 1963
rect 516 1937 668 1943
rect 964 1937 1020 1943
rect 1124 1937 1196 1943
rect 1220 1937 1324 1943
rect 1629 1937 1964 1943
rect 68 1917 332 1923
rect 436 1917 492 1923
rect 692 1917 764 1923
rect 772 1917 956 1923
rect 1012 1917 1116 1923
rect 1629 1923 1635 1937
rect 2132 1937 2188 1943
rect 2404 1937 2540 1943
rect 2644 1937 3132 1943
rect 3252 1937 4732 1943
rect 5140 1937 5644 1943
rect 5684 1937 5836 1943
rect 5860 1937 6092 1943
rect 6132 1937 6492 1943
rect 6500 1937 6604 1943
rect 1172 1917 1635 1923
rect 1652 1917 1708 1923
rect 1988 1917 2012 1923
rect 2020 1917 2124 1923
rect 2372 1917 2492 1923
rect 2612 1917 2812 1923
rect 2900 1917 3724 1923
rect 3860 1917 3964 1923
rect 3988 1917 4076 1923
rect 4116 1917 4140 1923
rect 4228 1917 4428 1923
rect 4436 1917 4588 1923
rect 4596 1917 4764 1923
rect 5012 1917 5148 1923
rect 5220 1917 5276 1923
rect 5284 1917 5532 1923
rect 5748 1917 5884 1923
rect 6020 1917 6076 1923
rect 6148 1917 6492 1923
rect 6740 1917 6860 1923
rect 6932 1917 6940 1923
rect 6964 1917 7100 1923
rect 116 1897 204 1903
rect 628 1897 716 1903
rect 980 1897 1004 1903
rect 1268 1897 1308 1903
rect 1348 1897 1372 1903
rect 1636 1897 1692 1903
rect 1796 1897 2076 1903
rect 2164 1897 2236 1903
rect 2260 1897 2284 1903
rect 2324 1897 2380 1903
rect 2740 1897 2764 1903
rect 2788 1897 2828 1903
rect 2900 1897 3020 1903
rect 3028 1897 3084 1903
rect 3092 1897 3180 1903
rect 3188 1897 3244 1903
rect 3252 1897 3308 1903
rect 3364 1897 3452 1903
rect 3556 1897 3612 1903
rect 3620 1897 3692 1903
rect 3700 1897 3868 1903
rect 3924 1897 4236 1903
rect 4244 1897 4364 1903
rect 4532 1897 4844 1903
rect 5316 1897 5516 1903
rect 5556 1897 5788 1903
rect 5924 1897 6044 1903
rect 6068 1897 6140 1903
rect 6148 1897 6179 1903
rect 20 1877 108 1883
rect 148 1877 300 1883
rect 500 1877 524 1883
rect 532 1877 684 1883
rect 724 1877 844 1883
rect 916 1877 1052 1883
rect 1092 1877 1324 1883
rect 1700 1877 1740 1883
rect 1876 1877 1900 1883
rect 1924 1877 1980 1883
rect 2260 1877 2268 1883
rect 2356 1877 2556 1883
rect 2916 1877 3036 1883
rect 3044 1877 3100 1883
rect 3108 1877 3196 1883
rect 3204 1877 3260 1883
rect 3268 1877 3324 1883
rect 3412 1877 3468 1883
rect 3492 1877 3676 1883
rect 3716 1877 3724 1883
rect 3748 1877 3804 1883
rect 3876 1877 3980 1883
rect 3988 1877 4044 1883
rect 4052 1877 4140 1883
rect 4276 1877 4300 1883
rect 4500 1877 4524 1883
rect 4532 1877 4604 1883
rect 4708 1877 4892 1883
rect 5028 1877 5132 1883
rect 5476 1877 5564 1883
rect 5572 1877 5619 1883
rect 148 1857 172 1863
rect 324 1857 428 1863
rect 644 1857 748 1863
rect 756 1857 860 1863
rect 932 1857 972 1863
rect 1044 1857 1068 1863
rect 1220 1857 1244 1863
rect 1364 1857 1964 1863
rect 1988 1857 2172 1863
rect 2196 1857 2428 1863
rect 2580 1857 2604 1863
rect 2836 1857 2876 1863
rect 3188 1857 3356 1863
rect 3380 1857 3692 1863
rect 3700 1857 3836 1863
rect 3940 1857 3980 1863
rect 4004 1857 4044 1863
rect 4148 1857 4188 1863
rect 4260 1857 4268 1863
rect 4308 1857 4524 1863
rect 4564 1857 4620 1863
rect 4724 1857 4748 1863
rect 5140 1857 5308 1863
rect 5460 1857 5580 1863
rect 5613 1863 5619 1877
rect 5636 1877 5772 1883
rect 5780 1877 6156 1883
rect 6173 1883 6179 1897
rect 6196 1897 6268 1903
rect 6292 1897 6892 1903
rect 6900 1897 6956 1903
rect 6996 1897 7068 1903
rect 6173 1877 6348 1883
rect 6356 1877 6396 1883
rect 6420 1877 6476 1883
rect 6484 1877 6508 1883
rect 6660 1877 6812 1883
rect 6852 1877 6892 1883
rect 6900 1877 7052 1883
rect 7124 1877 7244 1883
rect 5613 1857 5756 1863
rect 5764 1857 5964 1863
rect 5988 1857 6051 1863
rect 148 1837 156 1843
rect 260 1837 979 1843
rect 196 1817 396 1823
rect 452 1817 716 1823
rect 973 1823 979 1837
rect 996 1837 1004 1843
rect 1236 1837 1948 1843
rect 1972 1837 2060 1843
rect 2084 1837 2316 1843
rect 2356 1837 2396 1843
rect 2532 1837 2604 1843
rect 2628 1837 3036 1843
rect 3284 1837 3468 1843
rect 3508 1837 3628 1843
rect 3636 1837 3660 1843
rect 3684 1837 3788 1843
rect 3828 1837 4972 1843
rect 5124 1837 5228 1843
rect 5236 1837 5724 1843
rect 5764 1837 6028 1843
rect 6045 1843 6051 1857
rect 6100 1857 6108 1863
rect 6116 1857 6156 1863
rect 6164 1857 6204 1863
rect 6228 1857 6284 1863
rect 6324 1857 6508 1863
rect 6532 1857 6908 1863
rect 6916 1857 6956 1863
rect 7060 1857 7100 1863
rect 7188 1857 7219 1863
rect 6045 1837 6172 1843
rect 6285 1843 6291 1856
rect 6285 1837 6428 1843
rect 6468 1837 6956 1843
rect 7156 1837 7196 1843
rect 7213 1843 7219 1857
rect 7284 1857 7308 1863
rect 7213 1837 7276 1843
rect 7348 1837 7356 1843
rect 973 1817 1788 1823
rect 1860 1817 2092 1823
rect 2116 1817 2220 1823
rect 2244 1817 2844 1823
rect 3636 1817 4012 1823
rect 4308 1817 4364 1823
rect 5076 1817 5132 1823
rect 5140 1817 5388 1823
rect 5396 1817 5756 1823
rect 5780 1817 5868 1823
rect 6084 1817 6380 1823
rect 6420 1817 6428 1823
rect 6452 1817 6556 1823
rect 6740 1817 6748 1823
rect 6932 1817 6988 1823
rect 7188 1817 7372 1823
rect 2914 1814 2974 1816
rect 2914 1806 2915 1814
rect 2924 1806 2925 1814
rect 2963 1806 2964 1814
rect 2973 1806 2974 1814
rect 2914 1804 2974 1806
rect 5922 1814 5982 1816
rect 5922 1806 5923 1814
rect 5932 1806 5933 1814
rect 5971 1806 5972 1814
rect 5981 1806 5982 1814
rect 5922 1804 5982 1806
rect 212 1797 332 1803
rect 340 1797 1132 1803
rect 1300 1797 1356 1803
rect 1396 1797 1500 1803
rect 1524 1797 1836 1803
rect 1972 1797 2636 1803
rect 2692 1797 2844 1803
rect 3044 1797 3340 1803
rect 3396 1797 3500 1803
rect 3508 1797 3836 1803
rect 3853 1797 4844 1803
rect 580 1777 700 1783
rect 1124 1777 1292 1783
rect 1300 1777 1628 1783
rect 1652 1777 2284 1783
rect 2324 1777 2412 1783
rect 2468 1777 2668 1783
rect 2740 1777 2940 1783
rect 2948 1777 3388 1783
rect 3444 1777 3452 1783
rect 3508 1777 3532 1783
rect 3853 1783 3859 1797
rect 5252 1797 5660 1803
rect 6061 1797 6092 1803
rect 3652 1777 3859 1783
rect 3908 1777 4028 1783
rect 4244 1777 4300 1783
rect 4372 1777 4492 1783
rect 5588 1777 5596 1783
rect 5652 1777 5852 1783
rect 6061 1783 6067 1797
rect 6292 1797 6332 1803
rect 6596 1797 6652 1803
rect 7044 1797 7404 1803
rect 5908 1777 6067 1783
rect 6084 1777 6284 1783
rect 6324 1777 6764 1783
rect 7140 1777 7148 1783
rect 7188 1777 7324 1783
rect 7341 1764 7347 1776
rect 196 1757 236 1763
rect 276 1757 428 1763
rect 484 1757 1052 1763
rect 1092 1757 1148 1763
rect 1268 1757 1308 1763
rect 1348 1757 1356 1763
rect 1412 1757 1740 1763
rect 2004 1757 2492 1763
rect 2756 1757 2828 1763
rect 2836 1757 3372 1763
rect 3684 1757 3724 1763
rect 4068 1757 4140 1763
rect 4196 1757 4236 1763
rect 4244 1757 4460 1763
rect 4532 1757 4563 1763
rect 77 1737 172 1743
rect 77 1724 83 1737
rect 180 1737 476 1743
rect 580 1737 636 1743
rect 692 1737 700 1743
rect 916 1737 940 1743
rect 980 1737 1180 1743
rect 1188 1737 1548 1743
rect 1556 1737 1836 1743
rect 1844 1737 2252 1743
rect 2260 1737 2348 1743
rect 2628 1737 2796 1743
rect 2804 1737 3260 1743
rect 3284 1737 3356 1743
rect 3380 1737 3404 1743
rect 3476 1737 3507 1743
rect 68 1717 76 1723
rect 100 1717 204 1723
rect 228 1717 268 1723
rect 420 1717 451 1723
rect 68 1697 108 1703
rect 205 1703 211 1716
rect 205 1697 428 1703
rect 445 1703 451 1717
rect 548 1717 556 1723
rect 564 1717 620 1723
rect 628 1717 668 1723
rect 676 1717 780 1723
rect 1140 1717 1148 1723
rect 1156 1717 1516 1723
rect 1540 1717 1644 1723
rect 1684 1717 1788 1723
rect 1796 1717 1884 1723
rect 2004 1717 2108 1723
rect 2116 1717 2220 1723
rect 2276 1717 2284 1723
rect 2388 1717 2396 1723
rect 2404 1717 2604 1723
rect 2724 1717 2780 1723
rect 2852 1717 2892 1723
rect 3204 1717 3484 1723
rect 3501 1723 3507 1737
rect 3524 1737 3532 1743
rect 3556 1737 3900 1743
rect 3972 1737 4076 1743
rect 4084 1737 4124 1743
rect 4132 1737 4172 1743
rect 4180 1737 4316 1743
rect 4324 1737 4540 1743
rect 4557 1743 4563 1757
rect 4580 1757 4684 1763
rect 4932 1757 5068 1763
rect 5108 1757 5420 1763
rect 5428 1757 5532 1763
rect 5588 1757 5708 1763
rect 5748 1757 5820 1763
rect 5908 1757 6124 1763
rect 6132 1757 6204 1763
rect 6228 1757 6316 1763
rect 6324 1757 6364 1763
rect 6420 1757 6492 1763
rect 6548 1757 6636 1763
rect 6644 1757 6764 1763
rect 6868 1757 6924 1763
rect 7172 1757 7276 1763
rect 4557 1737 4620 1743
rect 4676 1737 4716 1743
rect 4724 1737 4780 1743
rect 4836 1737 4908 1743
rect 4948 1737 5036 1743
rect 5284 1737 5372 1743
rect 5492 1737 5772 1743
rect 5844 1737 5884 1743
rect 6068 1737 6172 1743
rect 6180 1737 6188 1743
rect 6260 1737 6300 1743
rect 6372 1737 6444 1743
rect 6564 1737 6604 1743
rect 6628 1737 6748 1743
rect 6765 1737 6812 1743
rect 3501 1717 3788 1723
rect 3812 1717 3932 1723
rect 4132 1717 4140 1723
rect 4212 1717 4460 1723
rect 4484 1717 4588 1723
rect 4596 1717 4604 1723
rect 4612 1717 4620 1723
rect 4788 1717 4988 1723
rect 5300 1717 5324 1723
rect 5348 1717 5452 1723
rect 5524 1717 6060 1723
rect 6132 1717 6220 1723
rect 6276 1717 6300 1723
rect 6308 1717 6476 1723
rect 6580 1717 6652 1723
rect 6660 1717 6700 1723
rect 6765 1723 6771 1737
rect 6980 1737 7027 1743
rect 6740 1717 6771 1723
rect 6836 1717 6892 1723
rect 6964 1717 6972 1723
rect 7021 1723 7027 1737
rect 7044 1737 7084 1743
rect 7021 1717 7036 1723
rect 7092 1717 7132 1723
rect 445 1697 828 1703
rect 1092 1697 1132 1703
rect 1997 1703 2003 1716
rect 1300 1697 2003 1703
rect 2068 1697 2188 1703
rect 2228 1697 2252 1703
rect 2404 1697 2460 1703
rect 2548 1697 2572 1703
rect 3156 1697 4508 1703
rect 4532 1697 4812 1703
rect 5636 1697 5676 1703
rect 5700 1697 6316 1703
rect 6452 1697 6588 1703
rect 6612 1697 6668 1703
rect 6676 1697 6828 1703
rect 7140 1697 7276 1703
rect 164 1677 236 1683
rect 324 1677 972 1683
rect 1508 1677 1692 1683
rect 1700 1677 1820 1683
rect 1828 1677 1868 1683
rect 1924 1677 2044 1683
rect 2164 1677 2172 1683
rect 2228 1677 2508 1683
rect 2884 1677 3324 1683
rect 3476 1677 3516 1683
rect 3572 1677 3612 1683
rect 3652 1677 3676 1683
rect 3796 1677 4620 1683
rect 4724 1677 4940 1683
rect 5412 1677 6284 1683
rect 6308 1677 6924 1683
rect 7060 1677 7164 1683
rect 36 1657 268 1663
rect 292 1657 460 1663
rect 948 1657 1580 1663
rect 1684 1657 1708 1663
rect 1764 1657 2124 1663
rect 2356 1657 2524 1663
rect 2676 1657 3788 1663
rect 4084 1657 4156 1663
rect 4212 1657 4380 1663
rect 4564 1657 4764 1663
rect 5204 1657 5292 1663
rect 5300 1657 5484 1663
rect 5508 1657 5692 1663
rect 5828 1657 5996 1663
rect 6324 1657 6684 1663
rect 6692 1657 7180 1663
rect 1492 1637 1660 1643
rect 1940 1637 1996 1643
rect 2372 1637 2572 1643
rect 2708 1637 3724 1643
rect 3796 1637 3996 1643
rect 4356 1637 4380 1643
rect 4404 1637 4444 1643
rect 4468 1637 4499 1643
rect 1524 1617 1612 1623
rect 1908 1617 2012 1623
rect 2708 1617 2764 1623
rect 2772 1617 2796 1623
rect 2804 1617 3020 1623
rect 3060 1617 3164 1623
rect 3252 1617 3324 1623
rect 3332 1617 3644 1623
rect 3652 1617 3708 1623
rect 3716 1617 3772 1623
rect 3780 1617 3884 1623
rect 3908 1617 4140 1623
rect 4493 1623 4499 1637
rect 4548 1637 4556 1643
rect 4692 1637 4924 1643
rect 4948 1637 5468 1643
rect 5572 1637 5644 1643
rect 6052 1637 6099 1643
rect 4493 1617 5420 1623
rect 5780 1617 5804 1623
rect 6004 1617 6076 1623
rect 6093 1623 6099 1637
rect 6148 1637 6444 1643
rect 6500 1637 7180 1643
rect 6093 1617 6572 1623
rect 6596 1617 6700 1623
rect 7156 1617 7180 1623
rect 1410 1614 1470 1616
rect 1410 1606 1411 1614
rect 1420 1606 1421 1614
rect 1459 1606 1460 1614
rect 1469 1606 1470 1614
rect 1410 1604 1470 1606
rect 4418 1614 4478 1616
rect 4418 1606 4419 1614
rect 4428 1606 4429 1614
rect 4467 1606 4468 1614
rect 4477 1606 4478 1614
rect 4418 1604 4478 1606
rect 2996 1597 3836 1603
rect 3956 1597 4204 1603
rect 4500 1597 4940 1603
rect 4980 1597 5324 1603
rect 5332 1597 5516 1603
rect 5524 1597 5868 1603
rect 5908 1597 6108 1603
rect 6628 1597 6700 1603
rect 6804 1597 7212 1603
rect 692 1577 780 1583
rect 788 1577 1068 1583
rect 1268 1577 1564 1583
rect 2740 1577 3900 1583
rect 3924 1577 3932 1583
rect 3988 1577 4268 1583
rect 4372 1577 4876 1583
rect 5284 1577 6204 1583
rect 6228 1577 6236 1583
rect 6484 1577 6508 1583
rect 6532 1577 6764 1583
rect 7028 1577 7068 1583
rect 7188 1577 7196 1583
rect 372 1557 2652 1563
rect 2660 1557 2940 1563
rect 2964 1557 3804 1563
rect 3812 1557 4108 1563
rect 4148 1557 4492 1563
rect 4516 1557 4700 1563
rect 5236 1557 5404 1563
rect 5428 1557 5900 1563
rect 6036 1557 6060 1563
rect 6100 1557 6188 1563
rect 6228 1557 6476 1563
rect 6484 1557 6652 1563
rect 6724 1557 7052 1563
rect 7284 1557 7308 1563
rect 420 1537 748 1543
rect 932 1537 972 1543
rect 1108 1537 1148 1543
rect 1364 1537 2620 1543
rect 2820 1537 2956 1543
rect 3060 1537 3980 1543
rect 4004 1537 4108 1543
rect 4116 1537 4332 1543
rect 4340 1537 4396 1543
rect 4404 1537 4652 1543
rect 4660 1537 4764 1543
rect 4772 1537 4828 1543
rect 4932 1537 5196 1543
rect 5268 1537 5996 1543
rect 6036 1537 6348 1543
rect 6356 1537 6476 1543
rect 6852 1537 6876 1543
rect 6948 1537 6956 1543
rect 6996 1537 7084 1543
rect 7204 1537 7228 1543
rect 7252 1537 7356 1543
rect 644 1517 684 1523
rect 852 1517 876 1523
rect 884 1517 924 1523
rect 1076 1517 1100 1523
rect 1796 1517 1836 1523
rect 2164 1517 2188 1523
rect 2356 1517 2444 1523
rect 3316 1517 3532 1523
rect 3556 1517 3820 1523
rect 3876 1517 4300 1523
rect 4308 1517 4588 1523
rect 4596 1517 4732 1523
rect 4868 1517 5004 1523
rect 5124 1517 5212 1523
rect 5220 1517 5388 1523
rect 5412 1517 5596 1523
rect 5620 1517 5900 1523
rect 5924 1517 5980 1523
rect 5988 1517 6044 1523
rect 6148 1517 6284 1523
rect 6404 1517 6563 1523
rect 6557 1504 6563 1517
rect 6868 1517 7340 1523
rect 292 1497 348 1503
rect 404 1497 540 1503
rect 548 1497 572 1503
rect 708 1497 764 1503
rect 772 1497 940 1503
rect 948 1497 1084 1503
rect 1316 1497 1548 1503
rect 1556 1497 1564 1503
rect 1604 1497 1724 1503
rect 1732 1497 1804 1503
rect 1876 1497 1932 1503
rect 1956 1497 2044 1503
rect 2052 1497 2252 1503
rect 2420 1497 2476 1503
rect 2484 1497 2572 1503
rect 2580 1497 2716 1503
rect 3204 1497 3228 1503
rect 3252 1497 3292 1503
rect 3428 1497 3436 1503
rect 3492 1497 3628 1503
rect 3732 1497 3740 1503
rect 3780 1497 3916 1503
rect 4020 1497 4124 1503
rect 4356 1497 4412 1503
rect 4420 1497 4636 1503
rect 4644 1497 4780 1503
rect 4788 1497 4844 1503
rect 5108 1497 5308 1503
rect 5332 1497 5372 1503
rect 5380 1497 5468 1503
rect 5476 1497 5532 1503
rect 5556 1497 6092 1503
rect 6132 1497 6332 1503
rect 6340 1497 6460 1503
rect 6564 1497 6764 1503
rect 6772 1497 6956 1503
rect 6996 1497 7036 1503
rect 7060 1497 7228 1503
rect 7236 1497 7244 1503
rect 173 1477 300 1483
rect 173 1464 179 1477
rect 500 1477 540 1483
rect 548 1477 572 1483
rect 820 1477 860 1483
rect 884 1477 908 1483
rect 980 1477 1036 1483
rect 1108 1477 1228 1483
rect 1332 1477 1500 1483
rect 1556 1477 1740 1483
rect 1876 1477 1900 1483
rect 1949 1483 1955 1496
rect 1908 1477 1955 1483
rect 2100 1477 2364 1483
rect 2372 1477 2412 1483
rect 2436 1477 2588 1483
rect 2612 1477 2668 1483
rect 2708 1477 2748 1483
rect 2756 1477 2812 1483
rect 3172 1477 3212 1483
rect 3220 1477 3292 1483
rect 3300 1477 3308 1483
rect 3316 1477 3356 1483
rect 3364 1477 3420 1483
rect 3444 1477 3548 1483
rect 3652 1477 3676 1483
rect 3716 1477 3788 1483
rect 3828 1477 4092 1483
rect 4212 1477 4236 1483
rect 4308 1477 4572 1483
rect 4596 1477 4620 1483
rect 4660 1477 4748 1483
rect 4884 1477 4892 1483
rect 4964 1477 5276 1483
rect 5309 1483 5315 1496
rect 5309 1477 5555 1483
rect 84 1457 172 1463
rect 196 1457 252 1463
rect 452 1457 492 1463
rect 500 1457 556 1463
rect 756 1457 828 1463
rect 852 1457 972 1463
rect 1076 1457 1260 1463
rect 1268 1457 1484 1463
rect 1540 1457 1612 1463
rect 1940 1457 2076 1463
rect 2244 1457 2316 1463
rect 2372 1457 2428 1463
rect 2452 1457 2556 1463
rect 2772 1457 3868 1463
rect 3924 1457 4044 1463
rect 4084 1457 4188 1463
rect 4244 1457 4508 1463
rect 4532 1457 4940 1463
rect 4957 1457 5260 1463
rect 116 1437 140 1443
rect 212 1437 316 1443
rect 436 1437 460 1443
rect 660 1437 1100 1443
rect 1108 1437 1164 1443
rect 1172 1437 1180 1443
rect 1220 1437 1260 1443
rect 1348 1437 1516 1443
rect 1524 1437 1580 1443
rect 1588 1437 1676 1443
rect 1716 1437 1756 1443
rect 2292 1437 2332 1443
rect 2532 1437 2540 1443
rect 3012 1437 3132 1443
rect 3348 1437 3388 1443
rect 3428 1437 3500 1443
rect 3508 1437 3580 1443
rect 3588 1437 3596 1443
rect 3604 1437 3660 1443
rect 3668 1437 3756 1443
rect 3860 1437 3980 1443
rect 4036 1437 4076 1443
rect 4957 1443 4963 1457
rect 5549 1463 5555 1477
rect 5572 1477 5692 1483
rect 5812 1477 5852 1483
rect 6196 1477 6364 1483
rect 6372 1477 6412 1483
rect 6452 1477 6492 1483
rect 6644 1477 6732 1483
rect 6788 1477 6876 1483
rect 6932 1477 7116 1483
rect 7172 1477 7244 1483
rect 7252 1477 7292 1483
rect 5549 1457 5612 1463
rect 6212 1457 6252 1463
rect 6276 1457 6284 1463
rect 6324 1457 6380 1463
rect 6452 1457 6460 1463
rect 6468 1457 6723 1463
rect 4100 1437 4963 1443
rect 5092 1437 5164 1443
rect 5172 1437 5308 1443
rect 5444 1437 5532 1443
rect 5876 1437 6140 1443
rect 6180 1437 6540 1443
rect 6596 1437 6684 1443
rect 6717 1443 6723 1457
rect 6740 1457 6988 1463
rect 7165 1463 7171 1476
rect 7092 1457 7171 1463
rect 6717 1437 6748 1443
rect 6756 1437 6780 1443
rect 6932 1437 7180 1443
rect 804 1417 2748 1423
rect 3124 1417 3148 1423
rect 3604 1417 3628 1423
rect 3684 1417 3708 1423
rect 3908 1417 4188 1423
rect 4260 1417 4300 1423
rect 4564 1417 4588 1423
rect 4804 1417 4972 1423
rect 4996 1417 5132 1423
rect 5268 1417 5420 1423
rect 5508 1417 5580 1423
rect 5652 1417 5692 1423
rect 6084 1417 6204 1423
rect 6244 1417 6348 1423
rect 6484 1417 6796 1423
rect 6804 1417 6860 1423
rect 6916 1417 7068 1423
rect 7076 1417 7148 1423
rect 2914 1414 2974 1416
rect 2914 1406 2915 1414
rect 2924 1406 2925 1414
rect 2963 1406 2964 1414
rect 2973 1406 2974 1414
rect 2914 1404 2974 1406
rect 5922 1414 5982 1416
rect 5922 1406 5923 1414
rect 5932 1406 5933 1414
rect 5971 1406 5972 1414
rect 5981 1406 5982 1414
rect 5922 1404 5982 1406
rect 564 1397 604 1403
rect 612 1397 668 1403
rect 676 1397 860 1403
rect 1236 1397 1260 1403
rect 1348 1397 1580 1403
rect 1604 1397 2012 1403
rect 2164 1397 2460 1403
rect 2468 1397 2492 1403
rect 2612 1397 2700 1403
rect 3092 1397 3196 1403
rect 3380 1397 3628 1403
rect 3636 1397 3772 1403
rect 3828 1397 5244 1403
rect 5540 1397 5715 1403
rect 5709 1384 5715 1397
rect 5732 1397 5884 1403
rect 6116 1397 6636 1403
rect 6676 1397 6764 1403
rect 6900 1397 7004 1403
rect 7108 1397 7340 1403
rect 372 1377 396 1383
rect 740 1377 1212 1383
rect 1300 1377 1660 1383
rect 1668 1377 2204 1383
rect 2253 1377 2364 1383
rect 2253 1364 2259 1377
rect 2644 1377 2716 1383
rect 2756 1377 3468 1383
rect 3485 1377 4044 1383
rect 84 1357 92 1363
rect 100 1357 140 1363
rect 148 1357 204 1363
rect 228 1357 300 1363
rect 324 1357 636 1363
rect 644 1357 700 1363
rect 1156 1357 1324 1363
rect 1412 1357 1596 1363
rect 1620 1357 1884 1363
rect 2036 1357 2076 1363
rect 2196 1357 2252 1363
rect 2356 1357 2556 1363
rect 2580 1357 2620 1363
rect 3108 1357 3148 1363
rect 3485 1363 3491 1377
rect 4244 1377 4444 1383
rect 4532 1377 4684 1383
rect 4820 1377 5212 1383
rect 5220 1377 5548 1383
rect 5716 1377 5772 1383
rect 5796 1377 6332 1383
rect 6356 1377 6396 1383
rect 6420 1377 6460 1383
rect 6500 1377 6732 1383
rect 3236 1357 3491 1363
rect 3524 1357 3628 1363
rect 3972 1357 3996 1363
rect 4020 1357 4076 1363
rect 4260 1357 4508 1363
rect 4756 1357 4812 1363
rect 4868 1357 4908 1363
rect 4932 1357 4940 1363
rect 4948 1357 5100 1363
rect 5284 1357 5644 1363
rect 5652 1357 5772 1363
rect 5956 1357 6060 1363
rect 6180 1357 6396 1363
rect 6436 1357 6604 1363
rect 6660 1357 6684 1363
rect 6772 1357 7116 1363
rect 148 1337 204 1343
rect 340 1337 508 1343
rect 756 1337 796 1343
rect 852 1337 908 1343
rect 1220 1337 1372 1343
rect 1380 1337 1804 1343
rect 1828 1337 1932 1343
rect 2132 1337 2140 1343
rect 2148 1337 2188 1343
rect 2292 1337 2508 1343
rect 2612 1337 2620 1343
rect 2676 1337 2764 1343
rect 2868 1337 2908 1343
rect 3060 1337 3100 1343
rect 3108 1337 3212 1343
rect 3236 1337 3324 1343
rect 3348 1337 3532 1343
rect 3572 1337 3788 1343
rect 3853 1337 3939 1343
rect 132 1317 220 1323
rect 244 1317 364 1323
rect 468 1317 492 1323
rect 900 1317 940 1323
rect 948 1317 1132 1323
rect 1268 1317 1756 1323
rect 2004 1317 2140 1323
rect 2228 1317 2380 1323
rect 2420 1317 2668 1323
rect 2756 1317 2796 1323
rect 3156 1317 3276 1323
rect 3332 1317 3452 1323
rect 3476 1317 3532 1323
rect 3540 1317 3612 1323
rect 3853 1323 3859 1337
rect 3732 1317 3859 1323
rect 3933 1323 3939 1337
rect 3956 1337 4012 1343
rect 4052 1337 6012 1343
rect 6052 1337 6220 1343
rect 6228 1337 6492 1343
rect 6500 1337 6812 1343
rect 6820 1337 6828 1343
rect 6852 1337 6924 1343
rect 7044 1337 7132 1343
rect 7140 1337 7308 1343
rect 3933 1317 3996 1323
rect 4004 1317 4140 1323
rect 4164 1317 4556 1323
rect 5092 1317 5164 1323
rect 5172 1317 5660 1323
rect 5684 1317 5788 1323
rect 5924 1317 6572 1323
rect 6580 1317 6796 1323
rect 6804 1317 6892 1323
rect 7156 1317 7228 1323
rect 548 1297 620 1303
rect 1012 1297 1372 1303
rect 1556 1297 1612 1303
rect 1636 1297 1868 1303
rect 1892 1297 2028 1303
rect 2052 1297 2172 1303
rect 2340 1297 2492 1303
rect 2516 1297 2524 1303
rect 2532 1297 2604 1303
rect 2820 1297 2860 1303
rect 2868 1297 2940 1303
rect 2948 1297 3260 1303
rect 3268 1297 3436 1303
rect 3572 1297 3660 1303
rect 3668 1297 3852 1303
rect 3876 1297 3916 1303
rect 3988 1297 4044 1303
rect 4084 1297 4268 1303
rect 4276 1297 4348 1303
rect 4372 1297 4652 1303
rect 4916 1297 4988 1303
rect 5300 1297 5692 1303
rect 6036 1297 6108 1303
rect 6164 1297 6252 1303
rect 6292 1297 6364 1303
rect 6596 1297 6604 1303
rect 6628 1297 6716 1303
rect 6900 1297 7036 1303
rect 68 1277 92 1283
rect 100 1277 284 1283
rect 372 1277 588 1283
rect 612 1277 668 1283
rect 836 1277 3244 1283
rect 3796 1277 3852 1283
rect 3972 1277 4060 1283
rect 4084 1277 4108 1283
rect 4228 1277 4604 1283
rect 4653 1283 4659 1296
rect 4653 1277 5100 1283
rect 5204 1277 6060 1283
rect 6100 1277 6108 1283
rect 6324 1277 6396 1283
rect 6532 1277 6748 1283
rect 6852 1277 6924 1283
rect 180 1257 300 1263
rect 980 1257 1004 1263
rect 1188 1257 2060 1263
rect 2356 1257 2364 1263
rect 2404 1257 2444 1263
rect 2452 1257 2588 1263
rect 2772 1257 2908 1263
rect 3220 1257 3244 1263
rect 3444 1257 3564 1263
rect 3748 1257 3836 1263
rect 3844 1257 4108 1263
rect 4548 1257 4620 1263
rect 4836 1257 5100 1263
rect 5108 1257 5116 1263
rect 5204 1257 5708 1263
rect 6036 1257 6044 1263
rect 6845 1263 6851 1276
rect 6468 1257 6851 1263
rect 1220 1237 1244 1243
rect 1284 1237 1324 1243
rect 1396 1237 2844 1243
rect 2852 1237 3244 1243
rect 3396 1237 3596 1243
rect 3604 1237 3980 1243
rect 4180 1237 4316 1243
rect 4436 1237 4540 1243
rect 4564 1237 5644 1243
rect 5668 1237 6188 1243
rect 6228 1237 6460 1243
rect 6580 1237 6860 1243
rect 804 1217 1212 1223
rect 1220 1217 1388 1223
rect 1492 1217 1612 1223
rect 1652 1217 1708 1223
rect 2068 1217 3020 1223
rect 3844 1217 3932 1223
rect 3956 1217 4348 1223
rect 4500 1217 6012 1223
rect 6100 1217 6172 1223
rect 6180 1217 6252 1223
rect 6564 1217 6908 1223
rect 1410 1214 1470 1216
rect 1410 1206 1411 1214
rect 1420 1206 1421 1214
rect 1459 1206 1460 1214
rect 1469 1206 1470 1214
rect 1410 1204 1470 1206
rect 4418 1214 4478 1216
rect 4418 1206 4419 1214
rect 4428 1206 4429 1214
rect 4467 1206 4468 1214
rect 4477 1206 4478 1214
rect 4418 1204 4478 1206
rect 1028 1197 1308 1203
rect 1364 1197 1388 1203
rect 1588 1197 1596 1203
rect 1604 1197 1948 1203
rect 1988 1197 2188 1203
rect 2196 1197 2396 1203
rect 2484 1197 2508 1203
rect 2628 1197 3500 1203
rect 3556 1197 4156 1203
rect 4516 1197 4924 1203
rect 5540 1197 5644 1203
rect 5748 1197 5884 1203
rect 6084 1197 6204 1203
rect 6212 1197 6268 1203
rect 6468 1197 6572 1203
rect 1012 1177 2236 1183
rect 2388 1177 2460 1183
rect 3860 1177 4012 1183
rect 4100 1177 4195 1183
rect 1060 1157 1532 1163
rect 1684 1157 1907 1163
rect 180 1137 364 1143
rect 740 1137 844 1143
rect 964 1137 972 1143
rect 1901 1143 1907 1157
rect 2244 1157 3052 1163
rect 3236 1157 3948 1163
rect 4164 1157 4172 1163
rect 4189 1163 4195 1177
rect 4292 1177 4428 1183
rect 4484 1177 4524 1183
rect 4676 1177 4796 1183
rect 5076 1177 5180 1183
rect 5188 1177 5452 1183
rect 5460 1177 5516 1183
rect 5572 1177 5596 1183
rect 5684 1177 5724 1183
rect 5828 1177 5980 1183
rect 6068 1177 6092 1183
rect 6436 1177 6796 1183
rect 4189 1157 4684 1163
rect 5476 1157 5788 1163
rect 5876 1157 6140 1163
rect 6164 1157 6556 1163
rect 7028 1157 7084 1163
rect 980 1137 1891 1143
rect 1901 1137 2572 1143
rect 1885 1124 1891 1137
rect 2580 1137 3100 1143
rect 3956 1137 3980 1143
rect 4004 1137 4092 1143
rect 4260 1137 4332 1143
rect 4356 1137 4492 1143
rect 4596 1137 4652 1143
rect 4660 1137 4732 1143
rect 4740 1137 4828 1143
rect 4845 1137 4860 1143
rect 196 1117 492 1123
rect 676 1117 956 1123
rect 964 1117 1020 1123
rect 1044 1117 1731 1123
rect -35 1097 12 1103
rect 228 1097 236 1103
rect 324 1097 364 1103
rect 404 1097 444 1103
rect 660 1097 684 1103
rect 916 1097 1068 1103
rect 1092 1097 1148 1103
rect 1156 1097 1260 1103
rect 1268 1097 1436 1103
rect 1572 1097 1660 1103
rect 1725 1103 1731 1117
rect 1748 1117 1772 1123
rect 1892 1117 2204 1123
rect 2301 1117 2460 1123
rect 2301 1103 2307 1117
rect 2868 1117 2892 1123
rect 3476 1117 3484 1123
rect 3700 1117 3884 1123
rect 3892 1117 4028 1123
rect 4356 1117 4364 1123
rect 4845 1123 4851 1137
rect 5028 1137 5132 1143
rect 5140 1137 5196 1143
rect 5204 1137 5244 1143
rect 5460 1137 5724 1143
rect 5732 1137 6188 1143
rect 6196 1137 6284 1143
rect 6292 1137 6380 1143
rect 6388 1137 6572 1143
rect 6980 1137 7116 1143
rect 4612 1117 4851 1123
rect 4868 1117 4908 1123
rect 5412 1117 5484 1123
rect 5508 1117 5580 1123
rect 5716 1117 5772 1123
rect 5924 1117 6364 1123
rect 6484 1117 6492 1123
rect 6500 1117 6540 1123
rect 6964 1117 6972 1123
rect 7060 1117 7244 1123
rect 7252 1117 7292 1123
rect 1725 1097 2307 1103
rect 2324 1097 2348 1103
rect 2356 1097 2556 1103
rect 2804 1097 2828 1103
rect 2916 1097 3212 1103
rect 3284 1097 3340 1103
rect 3476 1097 3532 1103
rect 3700 1097 3756 1103
rect 3940 1097 3964 1103
rect 3988 1097 4044 1103
rect 4276 1097 4332 1103
rect 4340 1097 4380 1103
rect 4452 1097 4508 1103
rect 4532 1097 4579 1103
rect 292 1077 428 1083
rect 868 1077 1036 1083
rect 1060 1077 1116 1083
rect 1124 1077 1228 1083
rect 1236 1077 1276 1083
rect 1364 1077 1372 1083
rect 1389 1077 1516 1083
rect 68 1057 268 1063
rect 276 1057 332 1063
rect 340 1057 396 1063
rect 404 1057 508 1063
rect 516 1057 540 1063
rect 564 1057 572 1063
rect 580 1057 636 1063
rect 644 1057 780 1063
rect 788 1057 988 1063
rect 996 1057 1084 1063
rect 1389 1063 1395 1077
rect 1732 1077 1836 1083
rect 1844 1077 1916 1083
rect 1924 1077 2092 1083
rect 2308 1077 2867 1083
rect 1252 1057 1395 1063
rect 1412 1057 1516 1063
rect 1524 1057 1676 1063
rect 1780 1057 1788 1063
rect 1796 1057 1852 1063
rect 1956 1057 2076 1063
rect 2132 1057 2332 1063
rect 2452 1057 2524 1063
rect 2532 1057 2540 1063
rect 2861 1063 2867 1077
rect 2884 1077 3180 1083
rect 3220 1077 3468 1083
rect 3540 1077 3548 1083
rect 3940 1077 4012 1083
rect 4020 1077 4060 1083
rect 4068 1077 4172 1083
rect 4196 1077 4284 1083
rect 4573 1083 4579 1097
rect 4596 1097 4652 1103
rect 4660 1097 4748 1103
rect 4756 1097 4844 1103
rect 4900 1097 5068 1103
rect 5332 1097 5340 1103
rect 5364 1097 5388 1103
rect 5597 1097 5660 1103
rect 4573 1077 4620 1083
rect 4708 1077 4844 1083
rect 5060 1077 5132 1083
rect 5332 1077 5436 1083
rect 5444 1077 5516 1083
rect 5597 1083 5603 1097
rect 5716 1097 5836 1103
rect 5892 1097 6172 1103
rect 6196 1097 6220 1103
rect 6532 1097 6684 1103
rect 6964 1097 7372 1103
rect 5524 1077 5603 1083
rect 5620 1077 5692 1083
rect 5764 1077 5852 1083
rect 5860 1077 6060 1083
rect 6100 1077 6140 1083
rect 6740 1077 6828 1083
rect 6836 1077 7100 1083
rect 7236 1077 7260 1083
rect 7316 1077 7324 1083
rect 2612 1057 2851 1063
rect 2861 1057 2908 1063
rect 164 1037 236 1043
rect 244 1037 284 1043
rect 324 1037 508 1043
rect 516 1037 828 1043
rect 980 1037 1164 1043
rect 1300 1037 1420 1043
rect 1524 1037 1612 1043
rect 1620 1037 1660 1043
rect 2436 1037 2620 1043
rect 2845 1043 2851 1057
rect 3460 1057 3500 1063
rect 4068 1057 4076 1063
rect 4148 1057 4524 1063
rect 4580 1057 4620 1063
rect 4788 1057 4828 1063
rect 5108 1057 5420 1063
rect 5540 1057 5724 1063
rect 5732 1057 6236 1063
rect 6244 1057 6300 1063
rect 6308 1057 6428 1063
rect 6708 1057 7020 1063
rect 7268 1057 7356 1063
rect 2845 1037 3244 1043
rect 3332 1037 3516 1043
rect 3876 1037 4188 1043
rect 4532 1037 4780 1043
rect 5220 1037 5372 1043
rect 5412 1037 5836 1043
rect 6036 1037 6108 1043
rect 6148 1037 6188 1043
rect 7316 1037 7356 1043
rect 372 1017 556 1023
rect 772 1017 796 1023
rect 804 1017 1052 1023
rect 1108 1017 1340 1023
rect 1540 1017 1676 1023
rect 1828 1017 1932 1023
rect 1940 1017 1996 1023
rect 2196 1017 2492 1023
rect 2548 1017 2876 1023
rect 2996 1017 3020 1023
rect 3028 1017 3580 1023
rect 3588 1017 3596 1023
rect 3780 1017 3868 1023
rect 4052 1017 5116 1023
rect 5524 1017 5676 1023
rect 6036 1017 6044 1023
rect 6084 1017 6140 1023
rect 6164 1017 6188 1023
rect 6212 1017 6332 1023
rect 6468 1017 6508 1023
rect 7300 1017 7372 1023
rect 2914 1014 2974 1016
rect 2914 1006 2915 1014
rect 2924 1006 2925 1014
rect 2963 1006 2964 1014
rect 2973 1006 2974 1014
rect 2914 1004 2974 1006
rect 5922 1014 5982 1016
rect 5922 1006 5923 1014
rect 5932 1006 5933 1014
rect 5971 1006 5972 1014
rect 5981 1006 5982 1014
rect 5922 1004 5982 1006
rect 228 997 748 1003
rect 804 997 876 1003
rect 1844 997 1900 1003
rect 1908 997 2028 1003
rect 2036 997 2076 1003
rect 2084 997 2204 1003
rect 2292 997 2348 1003
rect 2356 997 2636 1003
rect 2644 997 2892 1003
rect 2989 997 3500 1003
rect 132 977 156 983
rect 532 977 812 983
rect 820 977 876 983
rect 1284 977 2092 983
rect 2164 977 2188 983
rect 2228 977 2252 983
rect 2989 983 2995 997
rect 3652 997 3660 1003
rect 3732 997 3916 1003
rect 3924 997 4028 1003
rect 4116 997 4236 1003
rect 5396 997 5571 1003
rect 2820 977 2995 983
rect 3172 977 3196 983
rect 3380 977 3404 983
rect 3428 977 3484 983
rect 3812 977 3932 983
rect 4052 977 4092 983
rect 4132 977 4252 983
rect 4420 977 4668 983
rect 4692 977 4892 983
rect 5236 977 5548 983
rect 5565 983 5571 997
rect 6052 997 6124 1003
rect 6132 997 6252 1003
rect 5565 977 6236 983
rect 6404 977 6508 983
rect 6612 977 6764 983
rect 7172 977 7228 983
rect 7348 977 7372 983
rect 484 957 524 963
rect 532 957 588 963
rect 596 957 620 963
rect 628 957 652 963
rect 692 957 780 963
rect 788 957 860 963
rect 900 957 940 963
rect 964 957 1036 963
rect 1124 957 1228 963
rect 1316 957 1740 963
rect 1965 957 2380 963
rect 292 937 364 943
rect 372 937 652 943
rect 660 937 716 943
rect 964 937 1068 943
rect 1204 937 1276 943
rect 1965 943 1971 957
rect 2644 957 3116 963
rect 3124 957 3468 963
rect 3892 957 3916 963
rect 3924 957 4044 963
rect 4292 957 4643 963
rect 1300 937 1971 943
rect 1988 937 2540 943
rect 2852 937 3116 943
rect 3364 937 3372 943
rect 3460 937 3484 943
rect 3492 937 3516 943
rect 3524 937 3612 943
rect 3620 937 3692 943
rect 3700 937 3756 943
rect 3796 937 3820 943
rect 3828 937 3932 943
rect 3940 937 3964 943
rect 4324 937 4540 943
rect 4637 943 4643 957
rect 4660 957 4860 963
rect 4868 957 4924 963
rect 5108 957 5212 963
rect 5316 957 5452 963
rect 5476 957 5500 963
rect 5540 957 5580 963
rect 6196 957 6268 963
rect 6436 957 6620 963
rect 6676 957 6748 963
rect 6884 957 7116 963
rect 7252 957 7372 963
rect 4637 937 4748 943
rect 4868 937 4892 943
rect 5188 937 5276 943
rect 5492 937 5564 943
rect 5572 937 5660 943
rect 6132 937 6524 943
rect 6532 937 6684 943
rect 6788 937 6908 943
rect 6996 937 7340 943
rect 452 917 492 923
rect 580 917 668 923
rect 676 917 732 923
rect 932 917 1020 923
rect 1188 917 1260 923
rect 1444 917 1548 923
rect 1764 917 2060 923
rect 2100 917 2220 923
rect 2244 917 2300 923
rect 2308 917 2524 923
rect 2532 917 2668 923
rect 3204 917 3388 923
rect 3396 917 3676 923
rect 3684 917 4348 923
rect 4516 917 4748 923
rect 4788 917 4796 923
rect 4916 917 5020 923
rect 5172 917 5500 923
rect 5620 917 5708 923
rect 5780 917 5900 923
rect 6084 917 6156 923
rect 6484 917 6540 923
rect 6628 917 6812 923
rect 6900 917 6988 923
rect 6996 917 7052 923
rect 7060 917 7212 923
rect 7268 917 7308 923
rect -35 897 12 903
rect 340 897 364 903
rect 564 897 2604 903
rect 3764 897 3836 903
rect 3876 897 4012 903
rect 4100 897 4124 903
rect 4132 897 4316 903
rect 4580 897 4716 903
rect 4756 897 4764 903
rect 4996 897 5036 903
rect 5156 897 5315 903
rect 52 877 396 883
rect 868 877 1292 883
rect 1396 877 1612 883
rect 1828 877 1868 883
rect 2068 877 2108 883
rect 2132 877 2140 883
rect 2148 877 3036 883
rect 3044 877 3100 883
rect 3540 877 4540 883
rect 4596 877 4860 883
rect 5140 877 5180 883
rect 5309 883 5315 897
rect 5348 897 5484 903
rect 5524 897 5564 903
rect 5572 897 5804 903
rect 5908 897 6252 903
rect 6260 897 6412 903
rect 6900 897 6972 903
rect 6980 897 7004 903
rect 7252 897 7276 903
rect 5309 877 6076 883
rect 6516 877 6988 883
rect 7236 877 7276 883
rect 20 857 60 863
rect 468 857 492 863
rect 788 857 2060 863
rect 2164 857 2268 863
rect 2276 857 2412 863
rect 2436 857 2476 863
rect 2484 857 2572 863
rect 2628 857 3708 863
rect 3876 857 4364 863
rect 4612 857 4796 863
rect 4820 857 5379 863
rect 852 837 940 843
rect 1268 837 1276 843
rect 2061 843 2067 856
rect 2061 837 2652 843
rect 2692 837 3132 843
rect 3140 837 3564 843
rect 3732 837 4524 843
rect 4548 837 5356 843
rect 5373 843 5379 857
rect 5988 857 6332 863
rect 6580 857 6796 863
rect 5373 837 6364 843
rect 6676 837 6828 843
rect 6836 837 6924 843
rect 2004 817 2092 823
rect 2100 817 2172 823
rect 2180 817 2316 823
rect 2340 817 2748 823
rect 2900 817 3196 823
rect 3604 817 3644 823
rect 3652 817 3756 823
rect 3764 817 3868 823
rect 3988 817 4220 823
rect 4228 817 4252 823
rect 4500 817 6220 823
rect 6308 817 6940 823
rect 7268 817 7356 823
rect 1410 814 1470 816
rect 1410 806 1411 814
rect 1420 806 1421 814
rect 1459 806 1460 814
rect 1469 806 1470 814
rect 1410 804 1470 806
rect 4418 814 4478 816
rect 4418 806 4419 814
rect 4428 806 4429 814
rect 4467 806 4468 814
rect 4477 806 4478 814
rect 4418 804 4478 806
rect 932 797 1324 803
rect 2500 797 2524 803
rect 4708 797 4844 803
rect 5012 797 5196 803
rect 5268 797 5452 803
rect 5556 797 5628 803
rect 5636 797 5996 803
rect 6020 797 6060 803
rect 6244 797 6796 803
rect 7300 797 7356 803
rect 1172 777 1788 783
rect 1876 777 1964 783
rect 1972 777 2684 783
rect 2740 777 3020 783
rect 3028 777 3516 783
rect 4020 777 4156 783
rect 4404 777 4508 783
rect 4532 777 4812 783
rect 4884 777 4892 783
rect 5044 777 5116 783
rect 6260 777 6604 783
rect 6708 777 6844 783
rect 852 757 1020 763
rect 1044 757 1132 763
rect 1348 757 1516 763
rect 2260 757 2396 763
rect 2788 757 2924 763
rect 3508 757 4044 763
rect 4196 757 4236 763
rect 4276 757 4412 763
rect 5316 757 5548 763
rect 5828 757 6012 763
rect 6116 757 6700 763
rect 6964 757 7004 763
rect 324 737 540 743
rect 580 737 1340 743
rect 1636 737 1660 743
rect 1668 737 1948 743
rect 2308 737 2316 743
rect 2388 737 2572 743
rect 2580 737 2819 743
rect 116 717 156 723
rect 468 717 524 723
rect 820 717 876 723
rect 964 717 1036 723
rect 1172 717 1180 723
rect 1300 717 1324 723
rect 1540 717 1612 723
rect 1636 717 1772 723
rect 1956 717 1980 723
rect 2196 717 2236 723
rect 2420 717 2476 723
rect 2500 717 2572 723
rect 2628 717 2668 723
rect 2813 723 2819 737
rect 2836 737 2876 743
rect 2900 737 3020 743
rect 3988 737 4124 743
rect 4164 737 4332 743
rect 4724 737 4796 743
rect 4820 737 4956 743
rect 5332 737 5532 743
rect 5540 737 6268 743
rect 6292 737 6684 743
rect 6820 737 6860 743
rect 6916 737 6956 743
rect 7092 737 7228 743
rect 2813 717 2860 723
rect 2948 717 3068 723
rect 3812 717 3932 723
rect 4052 717 4076 723
rect 4228 717 4284 723
rect 4644 717 4748 723
rect 4788 717 4844 723
rect 4852 717 4940 723
rect 5812 717 6140 723
rect 6180 717 6284 723
rect 6292 717 6412 723
rect 6420 717 6476 723
rect 6724 717 6908 723
rect 372 697 412 703
rect 548 697 572 703
rect 580 697 668 703
rect 692 697 1228 703
rect 1252 697 1356 703
rect 1508 697 1692 703
rect 1700 697 1948 703
rect 1956 697 1996 703
rect 2132 697 2188 703
rect 2564 697 3155 703
rect 3149 684 3155 697
rect 3412 697 3484 703
rect 3492 697 3724 703
rect 3732 697 3804 703
rect 3860 697 3916 703
rect 3924 697 3964 703
rect 3972 697 4172 703
rect 4180 697 4252 703
rect 4740 697 4956 703
rect 5028 697 5164 703
rect 5252 697 5388 703
rect 5508 697 6028 703
rect 6036 697 6188 703
rect 6212 697 6284 703
rect 6564 697 6604 703
rect 6644 697 6700 703
rect 6740 697 6828 703
rect 6852 697 6956 703
rect 7076 697 7148 703
rect 7156 697 7212 703
rect 7220 697 7308 703
rect 68 677 140 683
rect 164 677 188 683
rect 292 677 460 683
rect 484 677 716 683
rect 916 677 940 683
rect 964 677 1004 683
rect 1060 677 1116 683
rect 1476 677 1548 683
rect 1604 677 1628 683
rect 1821 677 1852 683
rect 84 657 156 663
rect 308 657 364 663
rect 756 657 780 663
rect 788 657 796 663
rect 804 657 844 663
rect 852 657 972 663
rect 1044 657 1068 663
rect 1092 657 1148 663
rect 1348 657 1580 663
rect 1821 663 1827 677
rect 2228 677 2332 683
rect 2340 677 2844 683
rect 2852 677 3036 683
rect 3044 677 3084 683
rect 3156 677 3388 683
rect 3956 677 4108 683
rect 4116 677 4172 683
rect 4180 677 4220 683
rect 4228 677 4236 683
rect 4548 677 4700 683
rect 4788 677 4812 683
rect 4932 677 5084 683
rect 5460 677 5644 683
rect 5796 677 5836 683
rect 5940 677 6124 683
rect 6132 677 6476 683
rect 6548 677 6588 683
rect 6692 677 6780 683
rect 6804 677 6924 683
rect 6932 677 6956 683
rect 6964 677 7020 683
rect 1636 657 1827 663
rect 1844 657 2092 663
rect 2100 657 2268 663
rect 2292 657 2332 663
rect 2420 657 2524 663
rect 2548 657 2556 663
rect 2564 657 2636 663
rect 2900 657 3004 663
rect 3012 657 3052 663
rect 3908 657 3996 663
rect 4036 657 4044 663
rect 4052 657 4188 663
rect 4788 657 4844 663
rect 5044 657 5148 663
rect 5156 657 5260 663
rect 5748 657 5868 663
rect 6004 657 6252 663
rect 6260 657 6492 663
rect 6500 657 6748 663
rect 6756 657 6812 663
rect 6836 657 7116 663
rect 7204 657 7276 663
rect 84 637 252 643
rect 260 637 396 643
rect 404 637 476 643
rect 788 637 812 643
rect 1037 643 1043 656
rect 820 637 1043 643
rect 1716 637 1740 643
rect 2308 637 2732 643
rect 2916 637 3052 643
rect 3764 637 3836 643
rect 3997 643 4003 656
rect 3997 637 4156 643
rect 4212 637 5772 643
rect 5780 637 5884 643
rect 5901 637 6243 643
rect 244 617 1292 623
rect 1364 617 2204 623
rect 2484 617 2748 623
rect 3828 617 4067 623
rect 2914 614 2974 616
rect 2914 606 2915 614
rect 2924 606 2925 614
rect 2963 606 2964 614
rect 2973 606 2974 614
rect 2914 604 2974 606
rect 708 597 844 603
rect 1364 597 1516 603
rect 1636 597 1660 603
rect 1732 597 1788 603
rect 1844 597 1868 603
rect 1956 597 2284 603
rect 2292 597 2652 603
rect 3492 597 3788 603
rect 3908 597 4044 603
rect 4061 603 4067 617
rect 4157 623 4163 636
rect 4157 617 4204 623
rect 4820 617 4860 623
rect 4948 617 4972 623
rect 5124 617 5292 623
rect 5300 617 5372 623
rect 5588 617 5676 623
rect 5716 617 5740 623
rect 5901 623 5907 637
rect 5780 617 5907 623
rect 6237 623 6243 637
rect 6372 637 6540 643
rect 6564 637 6604 643
rect 6612 637 7308 643
rect 7316 637 7324 643
rect 6237 617 6444 623
rect 7108 617 7292 623
rect 5922 614 5982 616
rect 5922 606 5923 614
rect 5932 606 5933 614
rect 5971 606 5972 614
rect 5981 606 5982 614
rect 5922 604 5982 606
rect 4061 597 4492 603
rect 4660 597 4796 603
rect 5204 597 5212 603
rect 5412 597 5612 603
rect 5620 597 5900 603
rect 6884 597 6972 603
rect 6980 597 7148 603
rect 116 577 236 583
rect 996 577 1084 583
rect 1396 577 2140 583
rect 2452 577 2476 583
rect 2516 577 2924 583
rect 3620 577 3980 583
rect 4532 577 4716 583
rect 4820 577 4924 583
rect 5876 577 6124 583
rect 6164 577 6332 583
rect 6340 577 6348 583
rect 6452 577 6908 583
rect 6916 577 7052 583
rect 7124 577 7180 583
rect 36 557 60 563
rect 292 557 380 563
rect 564 557 684 563
rect 708 557 748 563
rect 868 557 908 563
rect 916 557 940 563
rect 948 557 1164 563
rect 1268 557 1484 563
rect 1540 557 1724 563
rect 1748 557 1836 563
rect 1844 557 1996 563
rect 2004 557 2028 563
rect 2036 557 2092 563
rect 2164 557 2188 563
rect 2228 557 2252 563
rect 2436 557 2476 563
rect 2596 557 2620 563
rect 2788 557 2835 563
rect 52 537 188 543
rect 196 537 348 543
rect 372 537 412 543
rect 420 537 508 543
rect 628 537 700 543
rect 756 537 1004 543
rect 1012 537 1292 543
rect 1316 537 1427 543
rect 52 517 268 523
rect 596 517 652 523
rect 660 517 876 523
rect 1044 517 1228 523
rect 1284 517 1404 523
rect 1421 523 1427 537
rect 1652 537 1708 543
rect 1780 537 1868 543
rect 2020 537 2108 543
rect 2116 537 2156 543
rect 2436 537 2492 543
rect 2660 537 2796 543
rect 2829 543 2835 557
rect 2852 557 2908 563
rect 2925 557 3036 563
rect 2925 543 2931 557
rect 3828 557 3868 563
rect 3924 557 3980 563
rect 4052 557 4076 563
rect 4756 557 4812 563
rect 4820 557 4876 563
rect 4884 557 4908 563
rect 4925 563 4931 576
rect 4925 557 5116 563
rect 5188 557 5212 563
rect 5220 557 5228 563
rect 5236 557 5308 563
rect 5316 557 5468 563
rect 5476 557 5788 563
rect 5956 557 6028 563
rect 6036 557 6140 563
rect 6788 557 6812 563
rect 6820 557 6924 563
rect 7156 557 7244 563
rect 2829 537 2931 543
rect 3028 537 3132 543
rect 3268 537 3420 543
rect 3588 537 3596 543
rect 3972 537 3980 543
rect 4660 537 4860 543
rect 5012 537 5404 543
rect 5412 537 5484 543
rect 6436 537 6460 543
rect 6468 537 6748 543
rect 6772 537 6844 543
rect 6852 537 6892 543
rect 1421 517 1596 523
rect 1828 517 1868 523
rect 1924 517 1964 523
rect 2068 517 2236 523
rect 2292 517 2364 523
rect 2372 517 2508 523
rect 2532 517 2716 523
rect 2756 517 2812 523
rect 3021 523 3027 536
rect 2884 517 3027 523
rect 3300 517 3468 523
rect 3748 517 3804 523
rect 3876 517 4012 523
rect 4020 517 4076 523
rect 4148 517 4284 523
rect 4372 517 4716 523
rect 4756 517 4812 523
rect 4868 517 4908 523
rect 5060 517 5196 523
rect 5268 517 5324 523
rect 5332 517 5388 523
rect 5476 517 5596 523
rect 5716 517 5788 523
rect 5812 517 5820 523
rect 6292 517 6380 523
rect 6532 517 6620 523
rect 6692 517 6860 523
rect 6868 517 7052 523
rect 7060 517 7244 523
rect 212 497 300 503
rect 340 497 380 503
rect 388 497 412 503
rect 676 497 716 503
rect 724 497 748 503
rect 852 497 876 503
rect 884 497 972 503
rect 1332 497 1356 503
rect 1588 497 1740 503
rect 2164 497 2188 503
rect 2404 497 2428 503
rect 2484 497 2540 503
rect 2644 497 3164 503
rect 3684 497 3932 503
rect 4020 497 4316 503
rect 4788 497 4844 503
rect 4964 497 5148 503
rect 5156 497 5212 503
rect 5812 497 6012 503
rect 6388 497 6428 503
rect 6436 497 6476 503
rect 6484 497 6492 503
rect 6500 497 6556 503
rect 6900 497 7036 503
rect 244 477 1052 483
rect 1060 477 1276 483
rect 1284 477 1340 483
rect 1508 477 1644 483
rect 2308 477 2348 483
rect 2452 477 2492 483
rect 2580 477 2908 483
rect 4180 477 4220 483
rect 4388 477 4908 483
rect 4916 477 4956 483
rect 5124 477 5436 483
rect 5444 477 5612 483
rect 5828 477 6060 483
rect 1476 457 1756 463
rect 4692 457 5020 463
rect 5220 457 5804 463
rect 4948 437 4972 443
rect 7012 437 7180 443
rect 2356 417 2636 423
rect 1410 414 1470 416
rect 1410 406 1411 414
rect 1420 406 1421 414
rect 1459 406 1460 414
rect 1469 406 1470 414
rect 1410 404 1470 406
rect 4418 414 4478 416
rect 4418 406 4419 414
rect 4428 406 4429 414
rect 4467 406 4468 414
rect 4477 406 4478 414
rect 4418 404 4478 406
rect 2468 397 2572 403
rect 2580 397 3052 403
rect 3060 397 3356 403
rect 3780 397 3852 403
rect 4132 397 4332 403
rect 372 377 780 383
rect 788 377 940 383
rect 1092 377 1548 383
rect 1876 377 1964 383
rect 2212 377 2316 383
rect 2516 377 2668 383
rect 3140 377 3164 383
rect 3508 377 3548 383
rect 3780 377 3852 383
rect 4100 377 4668 383
rect 6068 377 6204 383
rect 756 357 924 363
rect 941 357 988 363
rect 404 337 668 343
rect 941 343 947 357
rect 1348 357 1388 363
rect 1620 357 2028 363
rect 2276 357 2620 363
rect 2820 357 3116 363
rect 3124 357 3372 363
rect 3956 357 4092 363
rect 4164 357 4220 363
rect 4308 357 4476 363
rect 4836 357 4940 363
rect 4964 357 5276 363
rect 6404 357 7260 363
rect 852 337 947 343
rect 964 337 1116 343
rect 1268 337 1836 343
rect 1972 337 2131 343
rect 2125 324 2131 337
rect 2244 337 2380 343
rect 2388 337 2604 343
rect 2612 337 2636 343
rect 2644 337 2716 343
rect 3108 337 3340 343
rect 3892 337 4796 343
rect 4820 337 5180 343
rect 5188 337 5244 343
rect 5796 337 6012 343
rect 6372 337 6556 343
rect 6740 337 6828 343
rect 372 317 428 323
rect 580 317 684 323
rect 804 317 844 323
rect 900 317 956 323
rect 1012 317 1148 323
rect 1188 317 1404 323
rect 1636 317 1692 323
rect 1860 317 1932 323
rect 2148 317 2220 323
rect 2292 317 2364 323
rect 2916 317 3068 323
rect 3140 317 3212 323
rect 3668 317 3868 323
rect 3892 317 3996 323
rect 4004 317 4124 323
rect 4132 317 4172 323
rect 4180 317 4700 323
rect 4708 317 4908 323
rect 4916 317 5148 323
rect 5444 317 5596 323
rect 5604 317 5740 323
rect 5748 317 5788 323
rect 5796 317 5836 323
rect 5892 317 5996 323
rect 6196 317 6284 323
rect 6292 317 6332 323
rect 6356 317 6428 323
rect 6740 317 6844 323
rect 6980 317 7404 323
rect 116 297 236 303
rect 244 297 284 303
rect 356 297 572 303
rect 580 297 604 303
rect 772 297 780 303
rect 788 297 1020 303
rect 1172 297 1180 303
rect 1220 297 1260 303
rect 1348 297 1596 303
rect 1716 297 1804 303
rect 1812 297 2252 303
rect 2269 297 2364 303
rect 20 277 204 283
rect 404 277 460 283
rect 596 277 636 283
rect 660 277 700 283
rect 724 277 844 283
rect 868 277 908 283
rect 1236 277 1420 283
rect 1620 277 1836 283
rect 1860 277 1964 283
rect 1981 277 2172 283
rect 260 257 316 263
rect 324 257 524 263
rect 861 263 867 276
rect 532 257 867 263
rect 884 257 1132 263
rect 1140 257 1212 263
rect 1236 257 1596 263
rect 1604 257 1756 263
rect 1764 257 1964 263
rect 1981 263 1987 277
rect 2269 283 2275 297
rect 2516 297 2732 303
rect 2772 297 2844 303
rect 2852 297 2956 303
rect 3124 297 3148 303
rect 3156 297 3292 303
rect 3540 297 3932 303
rect 4052 297 4076 303
rect 4708 297 4748 303
rect 4820 297 4844 303
rect 5172 297 5644 303
rect 5668 297 6092 303
rect 6148 297 6220 303
rect 6228 297 6476 303
rect 6484 297 6572 303
rect 6804 297 7004 303
rect 7268 297 7372 303
rect 2196 277 2275 283
rect 2420 277 2540 283
rect 2692 277 2988 283
rect 2996 277 3148 283
rect 3156 277 3228 283
rect 3236 277 3276 283
rect 3412 277 4028 283
rect 4036 277 4044 283
rect 4212 277 4300 283
rect 4388 277 4540 283
rect 4628 277 4876 283
rect 4900 277 5068 283
rect 5108 277 5132 283
rect 5140 277 6700 283
rect 6708 277 7036 283
rect 7172 277 7196 283
rect 1972 257 1987 263
rect 2036 257 2092 263
rect 2164 257 2444 263
rect 2452 257 2476 263
rect 2484 257 2540 263
rect 2548 257 2700 263
rect 2708 257 2796 263
rect 2852 257 3068 263
rect 3236 257 3340 263
rect 3764 257 3788 263
rect 3812 257 3868 263
rect 3972 257 4044 263
rect 4068 257 4092 263
rect 4164 257 4332 263
rect 4388 257 4796 263
rect 4804 257 4924 263
rect 4980 257 5340 263
rect 5380 257 5436 263
rect 5492 257 5788 263
rect 5796 257 5884 263
rect 6004 257 6268 263
rect 6484 257 6876 263
rect 68 237 108 243
rect 132 237 188 243
rect 212 237 300 243
rect 436 237 652 243
rect 676 237 972 243
rect 980 237 1020 243
rect 1172 237 1292 243
rect 1540 237 1644 243
rect 1924 237 1980 243
rect 2100 237 2140 243
rect 2196 237 2412 243
rect 2420 237 2524 243
rect 2532 237 2588 243
rect 2596 237 2764 243
rect 3156 237 3180 243
rect 3844 237 3932 243
rect 4036 237 4588 243
rect 4724 237 4924 243
rect 4948 237 4956 243
rect 4996 237 5148 243
rect 5236 237 5740 243
rect 6269 243 6275 256
rect 6269 237 6540 243
rect 6548 237 6716 243
rect 468 217 627 223
rect 196 197 220 203
rect 340 197 604 203
rect 621 203 627 217
rect 644 217 812 223
rect 820 217 924 223
rect 1444 217 1660 223
rect 1668 217 1708 223
rect 1716 217 1884 223
rect 1892 217 2428 223
rect 2573 217 2876 223
rect 621 197 1084 203
rect 1332 197 1612 203
rect 1668 197 1868 203
rect 1876 197 1996 203
rect 2084 197 2236 203
rect 2573 203 2579 217
rect 4100 217 4172 223
rect 4804 217 5196 223
rect 5284 217 5308 223
rect 5316 217 5660 223
rect 6228 217 6412 223
rect 6420 217 6860 223
rect 2914 214 2974 216
rect 2914 206 2915 214
rect 2924 206 2925 214
rect 2963 206 2964 214
rect 2973 206 2974 214
rect 2914 204 2974 206
rect 5922 214 5982 216
rect 5922 206 5923 214
rect 5932 206 5933 214
rect 5971 206 5972 214
rect 5981 206 5982 214
rect 5922 204 5982 206
rect 2356 197 2579 203
rect 2596 197 2860 203
rect 3252 197 3852 203
rect 3940 197 4012 203
rect 4020 197 4172 203
rect 4180 197 4380 203
rect 4500 197 4819 203
rect 148 177 220 183
rect 420 177 508 183
rect 525 177 620 183
rect 164 157 332 163
rect 356 157 364 163
rect 525 163 531 177
rect 772 177 876 183
rect 916 177 1004 183
rect 1012 177 1036 183
rect 1316 177 1516 183
rect 1524 177 1532 183
rect 1540 177 1804 183
rect 1812 177 1996 183
rect 2116 177 2284 183
rect 2324 177 2492 183
rect 2724 177 2764 183
rect 2772 177 2812 183
rect 3044 177 3116 183
rect 3380 177 3820 183
rect 3860 177 3884 183
rect 3965 177 4076 183
rect 3965 164 3971 177
rect 4372 177 4620 183
rect 4749 177 4796 183
rect 4749 164 4755 177
rect 4813 183 4819 197
rect 4868 197 5468 203
rect 5652 197 5708 203
rect 5876 197 5900 203
rect 6628 197 6652 203
rect 6820 197 7388 203
rect 4813 177 4908 183
rect 4932 177 5356 183
rect 5668 177 5820 183
rect 6100 177 6284 183
rect 6292 177 6668 183
rect 6692 177 6732 183
rect 6932 177 7052 183
rect 516 157 531 163
rect 612 157 684 163
rect 692 157 732 163
rect 804 157 812 163
rect 1028 157 1228 163
rect 1636 157 1740 163
rect 1748 157 1820 163
rect 2020 157 2499 163
rect 20 137 44 143
rect 52 137 92 143
rect 100 137 572 143
rect 580 137 748 143
rect 756 137 860 143
rect 1124 137 1244 143
rect 1700 137 1852 143
rect 1860 137 1900 143
rect 1972 137 2028 143
rect 2045 137 2140 143
rect 84 117 124 123
rect 388 117 444 123
rect 452 117 540 123
rect 868 117 908 123
rect 1636 117 1676 123
rect 1748 117 1788 123
rect 1796 117 1868 123
rect 2045 123 2051 137
rect 2404 137 2476 143
rect 2493 143 2499 157
rect 2612 157 2668 163
rect 2740 157 3052 163
rect 3060 157 3340 163
rect 3668 157 3724 163
rect 3732 157 3916 163
rect 3924 157 3964 163
rect 4004 157 4044 163
rect 4260 157 4396 163
rect 4564 157 4748 163
rect 4772 157 5036 163
rect 5060 157 5708 163
rect 6388 157 6892 163
rect 6948 157 7084 163
rect 2493 137 2620 143
rect 2733 143 2739 156
rect 2644 137 2739 143
rect 2788 137 2908 143
rect 3012 137 3196 143
rect 3716 137 3836 143
rect 3844 137 4268 143
rect 4420 137 4572 143
rect 4644 137 4652 143
rect 4660 137 4700 143
rect 5012 137 5276 143
rect 5556 137 5692 143
rect 5732 137 5836 143
rect 6020 137 6060 143
rect 7044 137 7196 143
rect 7204 137 7340 143
rect 1988 117 2051 123
rect 2116 117 2284 123
rect 2292 117 2348 123
rect 2660 117 2684 123
rect 2772 117 2796 123
rect 3636 117 4508 123
rect 4516 117 4604 123
rect 4612 117 4652 123
rect 4692 117 5036 123
rect 5044 117 5116 123
rect 5124 117 5180 123
rect 5284 117 5340 123
rect 5412 117 5580 123
rect 5700 117 5788 123
rect 5860 117 6092 123
rect 7021 123 7027 136
rect 6852 117 7212 123
rect 36 97 204 103
rect 292 97 316 103
rect 452 97 492 103
rect 612 97 636 103
rect 1140 97 1548 103
rect 1556 97 1772 103
rect 1780 97 1932 103
rect 1940 97 2300 103
rect 4004 97 4060 103
rect 4596 97 4844 103
rect 6052 97 6156 103
rect 6644 97 6652 103
rect 6660 97 7068 103
rect 404 77 460 83
rect 1284 77 1468 83
rect 2292 77 2316 83
rect 4836 77 4860 83
rect 4868 77 4876 83
rect 4820 37 4892 43
rect 3476 17 3500 23
rect 3572 17 3596 23
rect 4068 17 4076 23
rect 1410 14 1470 16
rect 1410 6 1411 14
rect 1420 6 1421 14
rect 1459 6 1460 14
rect 1469 6 1470 14
rect 1410 4 1470 6
rect 4418 14 4478 16
rect 4418 6 4419 14
rect 4428 6 4429 14
rect 4467 6 4468 14
rect 4477 6 4478 14
rect 4418 4 4478 6
<< m4contact >>
rect 3436 5416 3444 5424
rect 3468 5416 3476 5424
rect 2916 5406 2923 5414
rect 2923 5406 2924 5414
rect 2928 5406 2933 5414
rect 2933 5406 2935 5414
rect 2935 5406 2936 5414
rect 2940 5406 2943 5414
rect 2943 5406 2945 5414
rect 2945 5406 2948 5414
rect 2952 5406 2953 5414
rect 2953 5406 2955 5414
rect 2955 5406 2960 5414
rect 2964 5406 2965 5414
rect 2965 5406 2972 5414
rect 5924 5406 5931 5414
rect 5931 5406 5932 5414
rect 5936 5406 5941 5414
rect 5941 5406 5943 5414
rect 5943 5406 5944 5414
rect 5948 5406 5951 5414
rect 5951 5406 5953 5414
rect 5953 5406 5956 5414
rect 5960 5406 5961 5414
rect 5961 5406 5963 5414
rect 5963 5406 5968 5414
rect 5972 5406 5973 5414
rect 5973 5406 5980 5414
rect 3564 5396 3572 5404
rect 5644 5396 5652 5404
rect 5324 5356 5332 5364
rect 5420 5356 5428 5364
rect 1612 5336 1620 5344
rect 1676 5296 1684 5304
rect 3212 5296 3220 5304
rect 4012 5296 4020 5304
rect 5324 5316 5332 5324
rect 5388 5316 5396 5324
rect 5356 5296 5364 5304
rect 5420 5296 5428 5304
rect 3436 5276 3444 5284
rect 5804 5256 5812 5264
rect 1412 5206 1419 5214
rect 1419 5206 1420 5214
rect 1424 5206 1429 5214
rect 1429 5206 1431 5214
rect 1431 5206 1432 5214
rect 1436 5206 1439 5214
rect 1439 5206 1441 5214
rect 1441 5206 1444 5214
rect 1448 5206 1449 5214
rect 1449 5206 1451 5214
rect 1451 5206 1456 5214
rect 1460 5206 1461 5214
rect 1461 5206 1468 5214
rect 4420 5206 4427 5214
rect 4427 5206 4428 5214
rect 4432 5206 4437 5214
rect 4437 5206 4439 5214
rect 4439 5206 4440 5214
rect 4444 5206 4447 5214
rect 4447 5206 4449 5214
rect 4449 5206 4452 5214
rect 4456 5206 4457 5214
rect 4457 5206 4459 5214
rect 4459 5206 4464 5214
rect 4468 5206 4469 5214
rect 4469 5206 4476 5214
rect 1900 5176 1908 5184
rect 2668 5176 2676 5184
rect 3436 5156 3444 5164
rect 5196 5156 5204 5164
rect 140 5136 148 5144
rect 4716 5136 4724 5144
rect 5740 5136 5748 5144
rect 4652 5116 4660 5124
rect 5708 5116 5716 5124
rect 204 5096 212 5104
rect 1324 5096 1332 5104
rect 1772 5096 1780 5104
rect 3532 5096 3540 5104
rect 5548 5096 5556 5104
rect 6188 5096 6196 5104
rect 6860 5096 6868 5104
rect 5164 5076 5172 5084
rect 5484 5076 5492 5084
rect 3436 5056 3444 5064
rect 7372 5076 7380 5084
rect 5740 5056 5748 5064
rect 972 5016 980 5024
rect 2572 5016 2580 5024
rect 7116 5036 7124 5044
rect 7308 5036 7316 5044
rect 5324 5016 5332 5024
rect 6380 5016 6388 5024
rect 2916 5006 2923 5014
rect 2923 5006 2924 5014
rect 2928 5006 2933 5014
rect 2933 5006 2935 5014
rect 2935 5006 2936 5014
rect 2940 5006 2943 5014
rect 2943 5006 2945 5014
rect 2945 5006 2948 5014
rect 2952 5006 2953 5014
rect 2953 5006 2955 5014
rect 2955 5006 2960 5014
rect 2964 5006 2965 5014
rect 2965 5006 2972 5014
rect 5924 5006 5931 5014
rect 5931 5006 5932 5014
rect 5936 5006 5941 5014
rect 5941 5006 5943 5014
rect 5943 5006 5944 5014
rect 5948 5006 5951 5014
rect 5951 5006 5953 5014
rect 5953 5006 5956 5014
rect 5960 5006 5961 5014
rect 5961 5006 5963 5014
rect 5963 5006 5968 5014
rect 5972 5006 5973 5014
rect 5973 5006 5980 5014
rect 4620 4996 4628 5004
rect 108 4976 116 4984
rect 2028 4976 2036 4984
rect 2412 4976 2420 4984
rect 5644 4976 5652 4984
rect 204 4956 212 4964
rect 332 4956 340 4964
rect 1276 4956 1284 4964
rect 1580 4956 1588 4964
rect 1900 4956 1908 4964
rect 3084 4956 3092 4964
rect 3788 4956 3796 4964
rect 5100 4956 5108 4964
rect 2252 4936 2260 4944
rect 2380 4936 2388 4944
rect 3404 4936 3412 4944
rect 4044 4936 4052 4944
rect 1260 4916 1268 4924
rect 1772 4916 1780 4924
rect 2060 4916 2068 4924
rect 1324 4896 1332 4904
rect 4620 4916 4628 4924
rect 4876 4916 4884 4924
rect 5388 4936 5396 4944
rect 5612 4936 5620 4944
rect 6956 4936 6964 4944
rect 5260 4916 5268 4924
rect 5708 4916 5716 4924
rect 3468 4896 3476 4904
rect 5100 4896 5108 4904
rect 6028 4896 6036 4904
rect 7116 4896 7124 4904
rect 1356 4856 1364 4864
rect 2028 4856 2036 4864
rect 2060 4856 2068 4864
rect 5004 4856 5012 4864
rect 972 4836 980 4844
rect 2412 4836 2420 4844
rect 3212 4836 3220 4844
rect 3468 4836 3476 4844
rect 3340 4816 3348 4824
rect 5356 4836 5364 4844
rect 5804 4836 5812 4844
rect 6188 4836 6196 4844
rect 5612 4816 5620 4824
rect 6060 4816 6068 4824
rect 1412 4806 1419 4814
rect 1419 4806 1420 4814
rect 1424 4806 1429 4814
rect 1429 4806 1431 4814
rect 1431 4806 1432 4814
rect 1436 4806 1439 4814
rect 1439 4806 1441 4814
rect 1441 4806 1444 4814
rect 1448 4806 1449 4814
rect 1449 4806 1451 4814
rect 1451 4806 1456 4814
rect 1460 4806 1461 4814
rect 1461 4806 1468 4814
rect 4420 4806 4427 4814
rect 4427 4806 4428 4814
rect 4432 4806 4437 4814
rect 4437 4806 4439 4814
rect 4439 4806 4440 4814
rect 4444 4806 4447 4814
rect 4447 4806 4449 4814
rect 4449 4806 4452 4814
rect 4456 4806 4457 4814
rect 4457 4806 4459 4814
rect 4459 4806 4464 4814
rect 4468 4806 4469 4814
rect 4469 4806 4476 4814
rect 3628 4796 3636 4804
rect 4524 4796 4532 4804
rect 2604 4776 2612 4784
rect 3500 4776 3508 4784
rect 1676 4756 1684 4764
rect 2572 4756 2580 4764
rect 5164 4776 5172 4784
rect 5484 4776 5492 4784
rect 4524 4756 4532 4764
rect 4780 4756 4788 4764
rect 1324 4736 1332 4744
rect 4108 4736 4116 4744
rect 5516 4736 5524 4744
rect 7148 4736 7156 4744
rect 844 4716 852 4724
rect 1964 4716 1972 4724
rect 5196 4716 5204 4724
rect 5548 4716 5556 4724
rect 1644 4696 1652 4704
rect 2284 4696 2292 4704
rect 3148 4696 3156 4704
rect 3596 4696 3604 4704
rect 4940 4696 4948 4704
rect 5868 4696 5876 4704
rect 6060 4696 6068 4704
rect 6572 4696 6580 4704
rect 140 4676 148 4684
rect 300 4676 308 4684
rect 4684 4676 4692 4684
rect 4716 4676 4724 4684
rect 5036 4676 5044 4684
rect 5804 4676 5812 4684
rect 5388 4656 5396 4664
rect 4524 4636 4532 4644
rect 4012 4616 4020 4624
rect 2916 4606 2923 4614
rect 2923 4606 2924 4614
rect 2928 4606 2933 4614
rect 2933 4606 2935 4614
rect 2935 4606 2936 4614
rect 2940 4606 2943 4614
rect 2943 4606 2945 4614
rect 2945 4606 2948 4614
rect 2952 4606 2953 4614
rect 2953 4606 2955 4614
rect 2955 4606 2960 4614
rect 2964 4606 2965 4614
rect 2965 4606 2972 4614
rect 5924 4606 5931 4614
rect 5931 4606 5932 4614
rect 5936 4606 5941 4614
rect 5941 4606 5943 4614
rect 5943 4606 5944 4614
rect 5948 4606 5951 4614
rect 5951 4606 5953 4614
rect 5953 4606 5956 4614
rect 5960 4606 5961 4614
rect 5961 4606 5963 4614
rect 5963 4606 5968 4614
rect 5972 4606 5973 4614
rect 5973 4606 5980 4614
rect 1964 4596 1972 4604
rect 1292 4576 1300 4584
rect 2380 4556 2388 4564
rect 3436 4596 3444 4604
rect 3788 4576 3796 4584
rect 4652 4576 4660 4584
rect 4780 4596 4788 4604
rect 7084 4596 7092 4604
rect 7276 4596 7284 4604
rect 4876 4576 4884 4584
rect 2764 4556 2772 4564
rect 3564 4556 3572 4564
rect 6028 4556 6036 4564
rect 6124 4556 6132 4564
rect 1708 4536 1716 4544
rect 2572 4536 2580 4544
rect 2604 4536 2612 4544
rect 3084 4536 3092 4544
rect 6316 4536 6324 4544
rect 6572 4536 6580 4544
rect 4588 4516 4596 4524
rect 5164 4516 5172 4524
rect 5612 4516 5620 4524
rect 6220 4516 6228 4524
rect 6924 4516 6932 4524
rect 7116 4516 7124 4524
rect 3468 4496 3476 4504
rect 3532 4496 3540 4504
rect 5356 4496 5364 4504
rect 6316 4496 6324 4504
rect 7212 4496 7220 4504
rect 1580 4476 1588 4484
rect 5260 4476 5268 4484
rect 6188 4476 6196 4484
rect 1644 4456 1652 4464
rect 5516 4456 5524 4464
rect 2796 4436 2804 4444
rect 3244 4436 3252 4444
rect 3500 4436 3508 4444
rect 4588 4436 4596 4444
rect 5004 4436 5012 4444
rect 5612 4436 5620 4444
rect 3276 4416 3284 4424
rect 3948 4416 3956 4424
rect 4524 4416 4532 4424
rect 5452 4416 5460 4424
rect 6188 4416 6196 4424
rect 1412 4406 1419 4414
rect 1419 4406 1420 4414
rect 1424 4406 1429 4414
rect 1429 4406 1431 4414
rect 1431 4406 1432 4414
rect 1436 4406 1439 4414
rect 1439 4406 1441 4414
rect 1441 4406 1444 4414
rect 1448 4406 1449 4414
rect 1449 4406 1451 4414
rect 1451 4406 1456 4414
rect 1460 4406 1461 4414
rect 1461 4406 1468 4414
rect 4420 4406 4427 4414
rect 4427 4406 4428 4414
rect 4432 4406 4437 4414
rect 4437 4406 4439 4414
rect 4439 4406 4440 4414
rect 4444 4406 4447 4414
rect 4447 4406 4449 4414
rect 4449 4406 4452 4414
rect 4456 4406 4457 4414
rect 4457 4406 4459 4414
rect 4459 4406 4464 4414
rect 4468 4406 4469 4414
rect 4469 4406 4476 4414
rect 3500 4396 3508 4404
rect 6316 4396 6324 4404
rect 780 4376 788 4384
rect 748 4356 756 4364
rect 4108 4356 4116 4364
rect 6124 4376 6132 4384
rect 6156 4376 6164 4384
rect 5132 4336 5140 4344
rect 5324 4336 5332 4344
rect 5388 4336 5396 4344
rect 6124 4336 6132 4344
rect 524 4316 532 4324
rect 876 4316 884 4324
rect 1228 4316 1236 4324
rect 7148 4316 7156 4324
rect 1068 4296 1076 4304
rect 1580 4296 1588 4304
rect 2124 4296 2132 4304
rect 5548 4296 5556 4304
rect 5580 4296 5588 4304
rect 5644 4296 5652 4304
rect 5772 4296 5780 4304
rect 5804 4296 5812 4304
rect 5868 4296 5876 4304
rect 6252 4296 6260 4304
rect 108 4276 116 4284
rect 908 4276 916 4284
rect 1708 4276 1716 4284
rect 1772 4276 1780 4284
rect 4876 4276 4884 4284
rect 6572 4276 6580 4284
rect 3724 4256 3732 4264
rect 5356 4256 5364 4264
rect 5740 4256 5748 4264
rect 1004 4236 1012 4244
rect 1772 4236 1780 4244
rect 2252 4236 2260 4244
rect 3340 4236 3348 4244
rect 3500 4236 3508 4244
rect 5644 4236 5652 4244
rect 3084 4216 3092 4224
rect 2916 4206 2923 4214
rect 2923 4206 2924 4214
rect 2928 4206 2933 4214
rect 2933 4206 2935 4214
rect 2935 4206 2936 4214
rect 2940 4206 2943 4214
rect 2943 4206 2945 4214
rect 2945 4206 2948 4214
rect 2952 4206 2953 4214
rect 2953 4206 2955 4214
rect 2955 4206 2960 4214
rect 2964 4206 2965 4214
rect 2965 4206 2972 4214
rect 5924 4206 5931 4214
rect 5931 4206 5932 4214
rect 5936 4206 5941 4214
rect 5941 4206 5943 4214
rect 5943 4206 5944 4214
rect 5948 4206 5951 4214
rect 5951 4206 5953 4214
rect 5953 4206 5956 4214
rect 5960 4206 5961 4214
rect 5961 4206 5963 4214
rect 5963 4206 5968 4214
rect 5972 4206 5973 4214
rect 5973 4206 5980 4214
rect 972 4196 980 4204
rect 2220 4196 2228 4204
rect 3372 4196 3380 4204
rect 3404 4196 3412 4204
rect 5580 4196 5588 4204
rect 5740 4196 5748 4204
rect 1036 4176 1044 4184
rect 5132 4176 5140 4184
rect 6284 4176 6292 4184
rect 6316 4176 6324 4184
rect 3468 4156 3476 4164
rect 4684 4156 4692 4164
rect 5836 4156 5844 4164
rect 6220 4156 6228 4164
rect 780 4136 788 4144
rect 1164 4136 1172 4144
rect 2572 4136 2580 4144
rect 3404 4136 3412 4144
rect 4364 4136 4372 4144
rect 5388 4136 5396 4144
rect 5644 4136 5652 4144
rect 5772 4136 5780 4144
rect 3628 4116 3636 4124
rect 3884 4116 3892 4124
rect 5868 4116 5876 4124
rect 6252 4116 6260 4124
rect 7244 4116 7252 4124
rect 1068 4096 1076 4104
rect 1164 4096 1172 4104
rect 2284 4096 2292 4104
rect 3244 4096 3252 4104
rect 5452 4096 5460 4104
rect 5676 4096 5684 4104
rect 5804 4096 5812 4104
rect 2412 4076 2420 4084
rect 2764 4076 2772 4084
rect 3084 4076 3092 4084
rect 5836 4076 5844 4084
rect 1324 4056 1332 4064
rect 1516 4056 1524 4064
rect 3116 4056 3124 4064
rect 2732 4036 2740 4044
rect 6444 4056 6452 4064
rect 7148 4056 7156 4064
rect 3148 4016 3156 4024
rect 6572 4016 6580 4024
rect 1412 4006 1419 4014
rect 1419 4006 1420 4014
rect 1424 4006 1429 4014
rect 1429 4006 1431 4014
rect 1431 4006 1432 4014
rect 1436 4006 1439 4014
rect 1439 4006 1441 4014
rect 1441 4006 1444 4014
rect 1448 4006 1449 4014
rect 1449 4006 1451 4014
rect 1451 4006 1456 4014
rect 1460 4006 1461 4014
rect 1461 4006 1468 4014
rect 4420 4006 4427 4014
rect 4427 4006 4428 4014
rect 4432 4006 4437 4014
rect 4437 4006 4439 4014
rect 4439 4006 4440 4014
rect 4444 4006 4447 4014
rect 4447 4006 4449 4014
rect 4449 4006 4452 4014
rect 4456 4006 4457 4014
rect 4457 4006 4459 4014
rect 4459 4006 4464 4014
rect 4468 4006 4469 4014
rect 4469 4006 4476 4014
rect 3468 3996 3476 4004
rect 6700 3996 6708 4004
rect 1356 3976 1364 3984
rect 1644 3976 1652 3984
rect 12 3956 20 3964
rect 3148 3976 3156 3984
rect 3308 3976 3316 3984
rect 3596 3976 3604 3984
rect 4588 3976 4596 3984
rect 6668 3976 6676 3984
rect 3276 3956 3284 3964
rect 5676 3956 5684 3964
rect 396 3936 404 3944
rect 1356 3936 1364 3944
rect 1676 3936 1684 3944
rect 172 3916 180 3924
rect 1036 3916 1044 3924
rect 1292 3916 1300 3924
rect 1708 3916 1716 3924
rect 4108 3916 4116 3924
rect 5772 3916 5780 3924
rect 908 3896 916 3904
rect 1548 3896 1556 3904
rect 1676 3896 1684 3904
rect 2476 3896 2484 3904
rect 2572 3896 2580 3904
rect 6892 3896 6900 3904
rect 2636 3876 2644 3884
rect 3884 3876 3892 3884
rect 5324 3876 5332 3884
rect 5772 3876 5780 3884
rect 6476 3876 6484 3884
rect 7020 3876 7028 3884
rect 972 3856 980 3864
rect 1004 3836 1012 3844
rect 5420 3856 5428 3864
rect 6252 3856 6260 3864
rect 6284 3856 6292 3864
rect 6060 3836 6068 3844
rect 6444 3836 6452 3844
rect 7244 3836 7252 3844
rect 812 3796 820 3804
rect 1292 3796 1300 3804
rect 4908 3816 4916 3824
rect 6956 3816 6964 3824
rect 7084 3816 7092 3824
rect 2916 3806 2923 3814
rect 2923 3806 2924 3814
rect 2928 3806 2933 3814
rect 2933 3806 2935 3814
rect 2935 3806 2936 3814
rect 2940 3806 2943 3814
rect 2943 3806 2945 3814
rect 2945 3806 2948 3814
rect 2952 3806 2953 3814
rect 2953 3806 2955 3814
rect 2955 3806 2960 3814
rect 2964 3806 2965 3814
rect 2965 3806 2972 3814
rect 5924 3806 5931 3814
rect 5931 3806 5932 3814
rect 5936 3806 5941 3814
rect 5941 3806 5943 3814
rect 5943 3806 5944 3814
rect 5948 3806 5951 3814
rect 5951 3806 5953 3814
rect 5953 3806 5956 3814
rect 5960 3806 5961 3814
rect 5961 3806 5963 3814
rect 5963 3806 5968 3814
rect 5972 3806 5973 3814
rect 5973 3806 5980 3814
rect 2508 3796 2516 3804
rect 3596 3796 3604 3804
rect 4204 3796 4212 3804
rect 4300 3796 4308 3804
rect 12 3756 20 3764
rect 876 3756 884 3764
rect 1036 3776 1044 3784
rect 3852 3776 3860 3784
rect 5612 3776 5620 3784
rect 6476 3776 6484 3784
rect 1356 3736 1364 3744
rect 2316 3736 2324 3744
rect 3692 3756 3700 3764
rect 4268 3756 4276 3764
rect 5324 3756 5332 3764
rect 7340 3776 7348 3784
rect 7244 3756 7252 3764
rect 5196 3736 5204 3744
rect 5388 3736 5396 3744
rect 5420 3736 5428 3744
rect 7084 3736 7092 3744
rect 172 3716 180 3724
rect 652 3716 660 3724
rect 812 3716 820 3724
rect 908 3716 916 3724
rect 2476 3716 2484 3724
rect 2636 3716 2644 3724
rect 3340 3716 3348 3724
rect 3852 3716 3860 3724
rect 4268 3716 4276 3724
rect 4940 3716 4948 3724
rect 5036 3716 5044 3724
rect 972 3676 980 3684
rect 4556 3696 4564 3704
rect 5100 3696 5108 3704
rect 6956 3716 6964 3724
rect 6444 3696 6452 3704
rect 6988 3696 6996 3704
rect 4908 3676 4916 3684
rect 6732 3676 6740 3684
rect 524 3656 532 3664
rect 5100 3656 5108 3664
rect 6092 3656 6100 3664
rect 844 3636 852 3644
rect 2668 3636 2676 3644
rect 3596 3636 3604 3644
rect 5740 3636 5748 3644
rect 6220 3636 6228 3644
rect 6700 3636 6708 3644
rect 6764 3636 6772 3644
rect 3724 3616 3732 3624
rect 1412 3606 1419 3614
rect 1419 3606 1420 3614
rect 1424 3606 1429 3614
rect 1429 3606 1431 3614
rect 1431 3606 1432 3614
rect 1436 3606 1439 3614
rect 1439 3606 1441 3614
rect 1441 3606 1444 3614
rect 1448 3606 1449 3614
rect 1449 3606 1451 3614
rect 1451 3606 1456 3614
rect 1460 3606 1461 3614
rect 1461 3606 1468 3614
rect 4420 3606 4427 3614
rect 4427 3606 4428 3614
rect 4432 3606 4437 3614
rect 4437 3606 4439 3614
rect 4439 3606 4440 3614
rect 4444 3606 4447 3614
rect 4447 3606 4449 3614
rect 4449 3606 4452 3614
rect 4456 3606 4457 3614
rect 4457 3606 4459 3614
rect 4459 3606 4464 3614
rect 4468 3606 4469 3614
rect 4469 3606 4476 3614
rect 1644 3596 1652 3604
rect 3372 3596 3380 3604
rect 6764 3596 6772 3604
rect 1932 3576 1940 3584
rect 3436 3576 3444 3584
rect 6572 3576 6580 3584
rect 7052 3576 7060 3584
rect 300 3536 308 3544
rect 1228 3536 1236 3544
rect 2572 3536 2580 3544
rect 3948 3536 3956 3544
rect 6028 3556 6036 3564
rect 6668 3556 6676 3564
rect 748 3516 756 3524
rect 1612 3516 1620 3524
rect 2476 3516 2484 3524
rect 3852 3516 3860 3524
rect 4108 3516 4116 3524
rect 6188 3516 6196 3524
rect 716 3496 724 3504
rect 876 3496 884 3504
rect 2060 3496 2068 3504
rect 2700 3496 2708 3504
rect 4300 3496 4308 3504
rect 4620 3496 4628 3504
rect 6060 3496 6068 3504
rect 6476 3496 6484 3504
rect 6892 3496 6900 3504
rect 332 3476 340 3484
rect 1708 3476 1716 3484
rect 1964 3476 1972 3484
rect 2316 3476 2324 3484
rect 2508 3476 2516 3484
rect 2732 3476 2740 3484
rect 3404 3476 3412 3484
rect 3884 3476 3892 3484
rect 6028 3476 6036 3484
rect 5164 3456 5172 3464
rect 1708 3436 1716 3444
rect 6028 3416 6036 3424
rect 2916 3406 2923 3414
rect 2923 3406 2924 3414
rect 2928 3406 2933 3414
rect 2933 3406 2935 3414
rect 2935 3406 2936 3414
rect 2940 3406 2943 3414
rect 2943 3406 2945 3414
rect 2945 3406 2948 3414
rect 2952 3406 2953 3414
rect 2953 3406 2955 3414
rect 2955 3406 2960 3414
rect 2964 3406 2965 3414
rect 2965 3406 2972 3414
rect 5924 3406 5931 3414
rect 5931 3406 5932 3414
rect 5936 3406 5941 3414
rect 5941 3406 5943 3414
rect 5943 3406 5944 3414
rect 5948 3406 5951 3414
rect 5951 3406 5953 3414
rect 5953 3406 5956 3414
rect 5960 3406 5961 3414
rect 5961 3406 5963 3414
rect 5963 3406 5968 3414
rect 5972 3406 5973 3414
rect 5973 3406 5980 3414
rect 876 3396 884 3404
rect 1900 3396 1908 3404
rect 6092 3396 6100 3404
rect 6188 3396 6196 3404
rect 780 3356 788 3364
rect 6124 3376 6132 3384
rect 2700 3356 2708 3364
rect 3116 3356 3124 3364
rect 3692 3356 3700 3364
rect 3724 3356 3732 3364
rect 5100 3356 5108 3364
rect 5452 3356 5460 3364
rect 7148 3356 7156 3364
rect 1356 3336 1364 3344
rect 6988 3336 6996 3344
rect 652 3316 660 3324
rect 1036 3316 1044 3324
rect 1868 3316 1876 3324
rect 4236 3316 4244 3324
rect 6636 3316 6644 3324
rect 7404 3316 7412 3324
rect 1612 3296 1620 3304
rect 1836 3296 1844 3304
rect 3116 3296 3124 3304
rect 3596 3296 3604 3304
rect 4076 3296 4084 3304
rect 4268 3296 4276 3304
rect 6156 3296 6164 3304
rect 5772 3276 5780 3284
rect 3340 3256 3348 3264
rect 3596 3256 3604 3264
rect 3660 3256 3668 3264
rect 7084 3256 7092 3264
rect 7212 3256 7220 3264
rect 5452 3236 5460 3244
rect 7276 3236 7284 3244
rect 1412 3206 1419 3214
rect 1419 3206 1420 3214
rect 1424 3206 1429 3214
rect 1429 3206 1431 3214
rect 1431 3206 1432 3214
rect 1436 3206 1439 3214
rect 1439 3206 1441 3214
rect 1441 3206 1444 3214
rect 1448 3206 1449 3214
rect 1449 3206 1451 3214
rect 1451 3206 1456 3214
rect 1460 3206 1461 3214
rect 1461 3206 1468 3214
rect 4420 3206 4427 3214
rect 4427 3206 4428 3214
rect 4432 3206 4437 3214
rect 4437 3206 4439 3214
rect 4439 3206 4440 3214
rect 4444 3206 4447 3214
rect 4447 3206 4449 3214
rect 4449 3206 4452 3214
rect 4456 3206 4457 3214
rect 4457 3206 4459 3214
rect 4459 3206 4464 3214
rect 4468 3206 4469 3214
rect 4469 3206 4476 3214
rect 2348 3196 2356 3204
rect 4140 3196 4148 3204
rect 5772 3196 5780 3204
rect 1548 3176 1556 3184
rect 1516 3156 1524 3164
rect 1932 3156 1940 3164
rect 2156 3156 2164 3164
rect 4588 3156 4596 3164
rect 5388 3156 5396 3164
rect 204 3116 212 3124
rect 396 3116 404 3124
rect 716 3116 724 3124
rect 748 3116 756 3124
rect 76 3096 84 3104
rect 364 3096 372 3104
rect 556 3096 564 3104
rect 4204 3136 4212 3144
rect 6988 3136 6996 3144
rect 1836 3116 1844 3124
rect 2572 3116 2580 3124
rect 6924 3116 6932 3124
rect 2412 3096 2420 3104
rect 4204 3096 4212 3104
rect 4716 3096 4724 3104
rect 5164 3096 5172 3104
rect 5452 3096 5460 3104
rect 6348 3096 6356 3104
rect 7052 3096 7060 3104
rect 588 3076 596 3084
rect 716 3076 724 3084
rect 780 3076 788 3084
rect 1036 3056 1044 3064
rect 4172 3076 4180 3084
rect 5196 3076 5204 3084
rect 6188 3076 6196 3084
rect 6284 3076 6292 3084
rect 6956 3076 6964 3084
rect 4204 3056 4212 3064
rect 4332 3056 4340 3064
rect 6924 3056 6932 3064
rect 908 3016 916 3024
rect 4300 3016 4308 3024
rect 6828 3016 6836 3024
rect 2916 3006 2923 3014
rect 2923 3006 2924 3014
rect 2928 3006 2933 3014
rect 2933 3006 2935 3014
rect 2935 3006 2936 3014
rect 2940 3006 2943 3014
rect 2943 3006 2945 3014
rect 2945 3006 2948 3014
rect 2952 3006 2953 3014
rect 2953 3006 2955 3014
rect 2955 3006 2960 3014
rect 2964 3006 2965 3014
rect 2965 3006 2972 3014
rect 5924 3006 5931 3014
rect 5931 3006 5932 3014
rect 5936 3006 5941 3014
rect 5941 3006 5943 3014
rect 5943 3006 5944 3014
rect 5948 3006 5951 3014
rect 5951 3006 5953 3014
rect 5953 3006 5956 3014
rect 5960 3006 5961 3014
rect 5961 3006 5963 3014
rect 5963 3006 5968 3014
rect 5972 3006 5973 3014
rect 5973 3006 5980 3014
rect 812 2996 820 3004
rect 2380 2996 2388 3004
rect 2700 2996 2708 3004
rect 4204 2996 4212 3004
rect 4364 2996 4372 3004
rect 3724 2976 3732 2984
rect 4012 2976 4020 2984
rect 7052 2976 7060 2984
rect 1676 2956 1684 2964
rect 3884 2956 3892 2964
rect 4556 2956 4564 2964
rect 6284 2956 6292 2964
rect 6476 2956 6484 2964
rect 6828 2956 6836 2964
rect 4332 2936 4340 2944
rect 6252 2936 6260 2944
rect 1036 2916 1044 2924
rect 1292 2916 1300 2924
rect 1868 2916 1876 2924
rect 2380 2916 2388 2924
rect 4172 2916 4180 2924
rect 4876 2916 4884 2924
rect 5548 2916 5556 2924
rect 5580 2916 5588 2924
rect 6220 2916 6228 2924
rect 7084 2916 7092 2924
rect 588 2896 596 2904
rect 1836 2896 1844 2904
rect 2060 2896 2068 2904
rect 3468 2896 3476 2904
rect 3820 2896 3828 2904
rect 3852 2896 3860 2904
rect 4204 2896 4212 2904
rect 4716 2896 4724 2904
rect 5836 2896 5844 2904
rect 1356 2876 1364 2884
rect 2476 2876 2484 2884
rect 3308 2876 3316 2884
rect 3372 2876 3380 2884
rect 4076 2876 4084 2884
rect 6796 2876 6804 2884
rect 364 2856 372 2864
rect 2444 2856 2452 2864
rect 4620 2856 4628 2864
rect 2156 2836 2164 2844
rect 3404 2836 3412 2844
rect 7180 2836 7188 2844
rect 1772 2816 1780 2824
rect 1804 2816 1812 2824
rect 2380 2816 2388 2824
rect 2636 2816 2644 2824
rect 1412 2806 1419 2814
rect 1419 2806 1420 2814
rect 1424 2806 1429 2814
rect 1429 2806 1431 2814
rect 1431 2806 1432 2814
rect 1436 2806 1439 2814
rect 1439 2806 1441 2814
rect 1441 2806 1444 2814
rect 1448 2806 1449 2814
rect 1449 2806 1451 2814
rect 1451 2806 1456 2814
rect 1460 2806 1461 2814
rect 1461 2806 1468 2814
rect 780 2776 788 2784
rect 876 2776 884 2784
rect 1516 2776 1524 2784
rect 1580 2776 1588 2784
rect 7404 2816 7412 2824
rect 4420 2806 4427 2814
rect 4427 2806 4428 2814
rect 4432 2806 4437 2814
rect 4437 2806 4439 2814
rect 4439 2806 4440 2814
rect 4444 2806 4447 2814
rect 4447 2806 4449 2814
rect 4449 2806 4452 2814
rect 4456 2806 4457 2814
rect 4457 2806 4459 2814
rect 4459 2806 4464 2814
rect 4468 2806 4469 2814
rect 4469 2806 4476 2814
rect 4268 2796 4276 2804
rect 4524 2796 4532 2804
rect 3756 2776 3764 2784
rect 1900 2756 1908 2764
rect 2700 2756 2708 2764
rect 3724 2756 3732 2764
rect 4684 2756 4692 2764
rect 7340 2756 7348 2764
rect 652 2736 660 2744
rect 748 2736 756 2744
rect 1708 2736 1716 2744
rect 2252 2736 2260 2744
rect 2700 2716 2708 2724
rect 3788 2736 3796 2744
rect 4076 2736 4084 2744
rect 4300 2736 4308 2744
rect 6764 2736 6772 2744
rect 3692 2716 3700 2724
rect 3724 2716 3732 2724
rect 7148 2716 7156 2724
rect 556 2696 564 2704
rect 1132 2696 1140 2704
rect 1164 2696 1172 2704
rect 1260 2696 1268 2704
rect 1580 2696 1588 2704
rect 1676 2696 1684 2704
rect 364 2676 372 2684
rect 2412 2676 2420 2684
rect 2476 2676 2484 2684
rect 2764 2676 2772 2684
rect 3916 2676 3924 2684
rect 4140 2696 4148 2704
rect 4204 2696 4212 2704
rect 4268 2676 4276 2684
rect 1228 2656 1236 2664
rect 1676 2656 1684 2664
rect 812 2636 820 2644
rect 844 2636 852 2644
rect 1900 2636 1908 2644
rect 1964 2656 1972 2664
rect 3724 2656 3732 2664
rect 3852 2656 3860 2664
rect 4012 2656 4020 2664
rect 4140 2656 4148 2664
rect 4588 2656 4596 2664
rect 7340 2696 7348 2704
rect 5740 2676 5748 2684
rect 6028 2676 6036 2684
rect 6284 2676 6292 2684
rect 5804 2656 5812 2664
rect 2220 2636 2228 2644
rect 2284 2636 2292 2644
rect 3436 2616 3444 2624
rect 4268 2616 4276 2624
rect 5836 2616 5844 2624
rect 2916 2606 2923 2614
rect 2923 2606 2924 2614
rect 2928 2606 2933 2614
rect 2933 2606 2935 2614
rect 2935 2606 2936 2614
rect 2940 2606 2943 2614
rect 2943 2606 2945 2614
rect 2945 2606 2948 2614
rect 2952 2606 2953 2614
rect 2953 2606 2955 2614
rect 2955 2606 2960 2614
rect 2964 2606 2965 2614
rect 2965 2606 2972 2614
rect 5924 2606 5931 2614
rect 5931 2606 5932 2614
rect 5936 2606 5941 2614
rect 5941 2606 5943 2614
rect 5943 2606 5944 2614
rect 5948 2606 5951 2614
rect 5951 2606 5953 2614
rect 5953 2606 5956 2614
rect 5960 2606 5961 2614
rect 5961 2606 5963 2614
rect 5963 2606 5968 2614
rect 5972 2606 5973 2614
rect 5973 2606 5980 2614
rect 3980 2596 3988 2604
rect 4108 2596 4116 2604
rect 4140 2596 4148 2604
rect 5228 2596 5236 2604
rect 3148 2576 3156 2584
rect 6732 2576 6740 2584
rect 460 2556 468 2564
rect 3788 2556 3796 2564
rect 4108 2556 4116 2564
rect 5804 2556 5812 2564
rect 2860 2536 2868 2544
rect 3916 2536 3924 2544
rect 4236 2536 4244 2544
rect 1996 2516 2004 2524
rect 2700 2516 2708 2524
rect 2796 2516 2804 2524
rect 3820 2516 3828 2524
rect 1324 2496 1332 2504
rect 2188 2496 2196 2504
rect 4076 2496 4084 2504
rect 4684 2536 4692 2544
rect 5548 2536 5556 2544
rect 4556 2516 4564 2524
rect 5228 2516 5236 2524
rect 5580 2516 5588 2524
rect 5644 2516 5652 2524
rect 6028 2516 6036 2524
rect 6444 2516 6452 2524
rect 6860 2516 6868 2524
rect 7276 2516 7284 2524
rect 4268 2496 4276 2504
rect 4588 2496 4596 2504
rect 4844 2496 4852 2504
rect 5612 2496 5620 2504
rect 780 2476 788 2484
rect 2124 2476 2132 2484
rect 2156 2476 2164 2484
rect 3692 2476 3700 2484
rect 4300 2476 4308 2484
rect 5644 2476 5652 2484
rect 5740 2476 5748 2484
rect 6956 2476 6964 2484
rect 1996 2456 2004 2464
rect 1580 2436 1588 2444
rect 2412 2436 2420 2444
rect 4108 2456 4116 2464
rect 4140 2456 4148 2464
rect 4364 2456 4372 2464
rect 4716 2456 4724 2464
rect 1004 2416 1012 2424
rect 1100 2416 1108 2424
rect 1324 2416 1332 2424
rect 1740 2416 1748 2424
rect 1772 2416 1780 2424
rect 1900 2416 1908 2424
rect 2604 2416 2612 2424
rect 5484 2436 5492 2444
rect 6700 2436 6708 2444
rect 4300 2416 4308 2424
rect 1412 2406 1419 2414
rect 1419 2406 1420 2414
rect 1424 2406 1429 2414
rect 1429 2406 1431 2414
rect 1431 2406 1432 2414
rect 1436 2406 1439 2414
rect 1439 2406 1441 2414
rect 1441 2406 1444 2414
rect 1448 2406 1449 2414
rect 1449 2406 1451 2414
rect 1451 2406 1456 2414
rect 1460 2406 1461 2414
rect 1461 2406 1468 2414
rect 4420 2406 4427 2414
rect 4427 2406 4428 2414
rect 4432 2406 4437 2414
rect 4437 2406 4439 2414
rect 4439 2406 4440 2414
rect 4444 2406 4447 2414
rect 4447 2406 4449 2414
rect 4449 2406 4452 2414
rect 4456 2406 4457 2414
rect 4457 2406 4459 2414
rect 4459 2406 4464 2414
rect 4468 2406 4469 2414
rect 4469 2406 4476 2414
rect 3916 2396 3924 2404
rect 4012 2396 4020 2404
rect 7212 2376 7220 2384
rect 172 2356 180 2364
rect 3468 2356 3476 2364
rect 3884 2356 3892 2364
rect 4044 2356 4052 2364
rect 4076 2356 4084 2364
rect 5484 2356 5492 2364
rect 5708 2356 5716 2364
rect 7372 2356 7380 2364
rect 780 2336 788 2344
rect 972 2336 980 2344
rect 1804 2336 1812 2344
rect 1964 2336 1972 2344
rect 3084 2336 3092 2344
rect 1996 2316 2004 2324
rect 2252 2316 2260 2324
rect 3116 2316 3124 2324
rect 684 2296 692 2304
rect 1260 2296 1268 2304
rect 1356 2296 1364 2304
rect 2092 2296 2100 2304
rect 2444 2296 2452 2304
rect 460 2276 468 2284
rect 1292 2276 1300 2284
rect 1836 2276 1844 2284
rect 2508 2276 2516 2284
rect 2764 2276 2772 2284
rect 3020 2276 3028 2284
rect 3532 2296 3540 2304
rect 3564 2296 3572 2304
rect 6764 2336 6772 2344
rect 4588 2316 4596 2324
rect 4748 2316 4756 2324
rect 5804 2316 5812 2324
rect 6284 2316 6292 2324
rect 3692 2276 3700 2284
rect 4588 2276 4596 2284
rect 4652 2276 4660 2284
rect 4716 2296 4724 2304
rect 5068 2296 5076 2304
rect 5612 2296 5620 2304
rect 4844 2276 4852 2284
rect 5644 2276 5652 2284
rect 6156 2296 6164 2304
rect 6572 2296 6580 2304
rect 7372 2296 7380 2304
rect 1164 2256 1172 2264
rect 2572 2256 2580 2264
rect 2604 2256 2612 2264
rect 2668 2256 2676 2264
rect 2700 2256 2708 2264
rect 3532 2256 3540 2264
rect 3948 2256 3956 2264
rect 2860 2236 2868 2244
rect 3660 2236 3668 2244
rect 3692 2236 3700 2244
rect 3756 2236 3764 2244
rect 3916 2236 3924 2244
rect 4076 2236 4084 2244
rect 1132 2216 1140 2224
rect 2732 2216 2740 2224
rect 4300 2216 4308 2224
rect 7404 2236 7412 2244
rect 5708 2216 5716 2224
rect 6220 2216 6228 2224
rect 2916 2206 2923 2214
rect 2923 2206 2924 2214
rect 2928 2206 2933 2214
rect 2933 2206 2935 2214
rect 2935 2206 2936 2214
rect 2940 2206 2943 2214
rect 2943 2206 2945 2214
rect 2945 2206 2948 2214
rect 2952 2206 2953 2214
rect 2953 2206 2955 2214
rect 2955 2206 2960 2214
rect 2964 2206 2965 2214
rect 2965 2206 2972 2214
rect 5924 2206 5931 2214
rect 5931 2206 5932 2214
rect 5936 2206 5941 2214
rect 5941 2206 5943 2214
rect 5943 2206 5944 2214
rect 5948 2206 5951 2214
rect 5951 2206 5953 2214
rect 5953 2206 5956 2214
rect 5960 2206 5961 2214
rect 5961 2206 5963 2214
rect 5963 2206 5968 2214
rect 5972 2206 5973 2214
rect 5973 2206 5980 2214
rect 7180 2216 7188 2224
rect 1196 2196 1204 2204
rect 2796 2196 2804 2204
rect 3692 2196 3700 2204
rect 4012 2196 4020 2204
rect 6668 2196 6676 2204
rect 6988 2196 6996 2204
rect 7052 2196 7060 2204
rect 2188 2176 2196 2184
rect 4268 2176 4276 2184
rect 4524 2176 4532 2184
rect 1356 2156 1364 2164
rect 2092 2156 2100 2164
rect 4076 2156 4084 2164
rect 4140 2156 4148 2164
rect 4972 2176 4980 2184
rect 6316 2176 6324 2184
rect 6924 2176 6932 2184
rect 5004 2156 5012 2164
rect 6220 2156 6228 2164
rect 1324 2136 1332 2144
rect 1964 2136 1972 2144
rect 2572 2136 2580 2144
rect 3852 2136 3860 2144
rect 4364 2136 4372 2144
rect 6348 2136 6356 2144
rect 6956 2136 6964 2144
rect 524 2116 532 2124
rect 652 2116 660 2124
rect 1228 2096 1236 2104
rect 1868 2096 1876 2104
rect 2828 2116 2836 2124
rect 3020 2116 3028 2124
rect 3244 2116 3252 2124
rect 3628 2116 3636 2124
rect 3724 2116 3732 2124
rect 3788 2116 3796 2124
rect 4012 2116 4020 2124
rect 4268 2116 4276 2124
rect 4652 2116 4660 2124
rect 4716 2116 4724 2124
rect 6860 2116 6868 2124
rect 7116 2116 7124 2124
rect 2252 2096 2260 2104
rect 2540 2096 2548 2104
rect 2636 2096 2644 2104
rect 2732 2096 2740 2104
rect 2796 2096 2804 2104
rect 3116 2096 3124 2104
rect 4300 2096 4308 2104
rect 172 2056 180 2064
rect 4076 2076 4084 2084
rect 4684 2076 4692 2084
rect 6156 2076 6164 2084
rect 1260 2056 1268 2064
rect 2316 2056 2324 2064
rect 2380 2056 2388 2064
rect 2508 2056 2516 2064
rect 2732 2056 2740 2064
rect 2764 2056 2772 2064
rect 716 2036 724 2044
rect 1228 2036 1236 2044
rect 3372 2036 3380 2044
rect 3596 2036 3604 2044
rect 6156 2036 6164 2044
rect 6828 2036 6836 2044
rect 7180 2036 7188 2044
rect 1868 2016 1876 2024
rect 3788 2016 3796 2024
rect 5100 2016 5108 2024
rect 6284 2016 6292 2024
rect 1412 2006 1419 2014
rect 1419 2006 1420 2014
rect 1424 2006 1429 2014
rect 1429 2006 1431 2014
rect 1431 2006 1432 2014
rect 1436 2006 1439 2014
rect 1439 2006 1441 2014
rect 1441 2006 1444 2014
rect 1448 2006 1449 2014
rect 1449 2006 1451 2014
rect 1451 2006 1456 2014
rect 1460 2006 1461 2014
rect 1461 2006 1468 2014
rect 4420 2006 4427 2014
rect 4427 2006 4428 2014
rect 4432 2006 4437 2014
rect 4437 2006 4439 2014
rect 4439 2006 4440 2014
rect 4444 2006 4447 2014
rect 4447 2006 4449 2014
rect 4449 2006 4452 2014
rect 4456 2006 4457 2014
rect 4457 2006 4459 2014
rect 4459 2006 4464 2014
rect 4468 2006 4469 2014
rect 4469 2006 4476 2014
rect 1196 1996 1204 2004
rect 2316 1996 2324 2004
rect 7116 1996 7124 2004
rect 5580 1976 5588 1984
rect 780 1956 788 1964
rect 3724 1956 3732 1964
rect 6412 1956 6420 1964
rect 2188 1936 2196 1944
rect 2636 1936 2644 1944
rect 1708 1916 1716 1924
rect 3724 1916 3732 1924
rect 3980 1916 3988 1924
rect 4140 1916 4148 1924
rect 6924 1916 6932 1924
rect 2380 1896 2388 1904
rect 4236 1896 4244 1904
rect 6060 1896 6068 1904
rect 524 1876 532 1884
rect 2252 1876 2260 1884
rect 2348 1876 2356 1884
rect 3724 1876 3732 1884
rect 4204 1876 4212 1884
rect 4300 1876 4308 1884
rect 4524 1876 4532 1884
rect 2188 1856 2196 1864
rect 2572 1856 2580 1864
rect 2604 1856 2612 1864
rect 2828 1856 2836 1864
rect 3372 1856 3380 1864
rect 3692 1856 3700 1864
rect 4076 1856 4084 1864
rect 4140 1856 4148 1864
rect 4268 1856 4276 1864
rect 5772 1876 5780 1884
rect 6156 1876 6164 1884
rect 6892 1896 6900 1904
rect 6988 1896 6996 1904
rect 7308 1896 7316 1904
rect 6572 1876 6580 1884
rect 7052 1876 7060 1884
rect 7116 1876 7124 1884
rect 140 1836 148 1844
rect 1004 1836 1012 1844
rect 1964 1836 1972 1844
rect 2316 1836 2324 1844
rect 2348 1836 2356 1844
rect 3500 1836 3508 1844
rect 4972 1836 4980 1844
rect 6028 1836 6036 1844
rect 6092 1856 6100 1864
rect 6316 1856 6324 1864
rect 6956 1836 6964 1844
rect 7308 1856 7316 1864
rect 7340 1836 7348 1844
rect 2220 1816 2228 1824
rect 4300 1816 4308 1824
rect 5068 1816 5076 1824
rect 5132 1816 5140 1824
rect 6412 1816 6420 1824
rect 6444 1816 6452 1824
rect 6668 1816 6676 1824
rect 6732 1816 6740 1824
rect 2916 1806 2923 1814
rect 2923 1806 2924 1814
rect 2928 1806 2933 1814
rect 2933 1806 2935 1814
rect 2935 1806 2936 1814
rect 2940 1806 2943 1814
rect 2943 1806 2945 1814
rect 2945 1806 2948 1814
rect 2952 1806 2953 1814
rect 2953 1806 2955 1814
rect 2955 1806 2960 1814
rect 2964 1806 2965 1814
rect 2965 1806 2972 1814
rect 5924 1806 5931 1814
rect 5931 1806 5932 1814
rect 5936 1806 5941 1814
rect 5941 1806 5943 1814
rect 5943 1806 5944 1814
rect 5948 1806 5951 1814
rect 5951 1806 5953 1814
rect 5953 1806 5956 1814
rect 5960 1806 5961 1814
rect 5961 1806 5963 1814
rect 5963 1806 5968 1814
rect 5972 1806 5973 1814
rect 5973 1806 5980 1814
rect 1132 1796 1140 1804
rect 2636 1796 2644 1804
rect 940 1776 948 1784
rect 1292 1776 1300 1784
rect 1644 1776 1652 1784
rect 2316 1776 2324 1784
rect 3436 1776 3444 1784
rect 3532 1776 3540 1784
rect 4300 1776 4308 1784
rect 5580 1776 5588 1784
rect 6284 1776 6292 1784
rect 6316 1776 6324 1784
rect 7148 1776 7156 1784
rect 7180 1776 7188 1784
rect 268 1756 276 1764
rect 1324 1756 1332 1764
rect 1356 1756 1364 1764
rect 3372 1756 3380 1764
rect 3916 1756 3924 1764
rect 4012 1756 4020 1764
rect 684 1736 692 1744
rect 972 1736 980 1744
rect 1836 1736 1844 1744
rect 2572 1736 2580 1744
rect 3404 1736 3412 1744
rect 76 1716 84 1724
rect 204 1716 212 1724
rect 268 1716 276 1724
rect 1004 1716 1012 1724
rect 1132 1716 1140 1724
rect 1644 1716 1652 1724
rect 1676 1716 1684 1724
rect 1964 1716 1972 1724
rect 1996 1716 2004 1724
rect 2284 1716 2292 1724
rect 2380 1716 2388 1724
rect 3532 1736 3540 1744
rect 5100 1756 5108 1764
rect 5548 1756 5556 1764
rect 6764 1756 6772 1764
rect 7340 1756 7348 1764
rect 6188 1736 6196 1744
rect 6444 1736 6452 1744
rect 3788 1716 3796 1724
rect 4140 1716 4148 1724
rect 4204 1716 4212 1724
rect 4588 1716 4596 1724
rect 6124 1716 6132 1724
rect 6572 1716 6580 1724
rect 6828 1716 6836 1724
rect 6956 1716 6964 1724
rect 7148 1736 7156 1744
rect 2252 1696 2260 1704
rect 4812 1696 4820 1704
rect 6316 1696 6324 1704
rect 6604 1696 6612 1704
rect 972 1676 980 1684
rect 1356 1676 1364 1684
rect 2156 1676 2164 1684
rect 2220 1676 2228 1684
rect 3564 1676 3572 1684
rect 3692 1676 3700 1684
rect 3788 1676 3796 1684
rect 2668 1656 2676 1664
rect 4076 1656 4084 1664
rect 5196 1656 5204 1664
rect 1708 1636 1716 1644
rect 2572 1636 2580 1644
rect 2700 1636 2708 1644
rect 3788 1636 3796 1644
rect 1516 1616 1524 1624
rect 1612 1616 1620 1624
rect 3020 1616 3028 1624
rect 3052 1616 3060 1624
rect 4140 1616 4148 1624
rect 4556 1636 4564 1644
rect 4940 1636 4948 1644
rect 5772 1616 5780 1624
rect 7180 1636 7188 1644
rect 1412 1606 1419 1614
rect 1419 1606 1420 1614
rect 1424 1606 1429 1614
rect 1429 1606 1431 1614
rect 1431 1606 1432 1614
rect 1436 1606 1439 1614
rect 1439 1606 1441 1614
rect 1441 1606 1444 1614
rect 1448 1606 1449 1614
rect 1449 1606 1451 1614
rect 1451 1606 1456 1614
rect 1460 1606 1461 1614
rect 1461 1606 1468 1614
rect 4420 1606 4427 1614
rect 4427 1606 4428 1614
rect 4432 1606 4437 1614
rect 4437 1606 4439 1614
rect 4439 1606 4440 1614
rect 4444 1606 4447 1614
rect 4447 1606 4449 1614
rect 4449 1606 4452 1614
rect 4456 1606 4457 1614
rect 4457 1606 4459 1614
rect 4459 1606 4464 1614
rect 4468 1606 4469 1614
rect 4469 1606 4476 1614
rect 4204 1596 4212 1604
rect 4940 1596 4948 1604
rect 5324 1596 5332 1604
rect 6700 1596 6708 1604
rect 6796 1596 6804 1604
rect 2732 1576 2740 1584
rect 3916 1576 3924 1584
rect 3948 1576 3956 1584
rect 3980 1576 3988 1584
rect 6220 1576 6228 1584
rect 6476 1576 6484 1584
rect 7180 1576 7188 1584
rect 4140 1556 4148 1564
rect 6028 1556 6036 1564
rect 7308 1556 7316 1564
rect 972 1536 980 1544
rect 1356 1536 1364 1544
rect 3980 1536 3988 1544
rect 5260 1536 5268 1544
rect 6476 1536 6484 1544
rect 6956 1536 6964 1544
rect 7244 1536 7252 1544
rect 1100 1516 1108 1524
rect 2188 1516 2196 1524
rect 3820 1516 3828 1524
rect 5612 1516 5620 1524
rect 6860 1516 6868 1524
rect 940 1496 948 1504
rect 1548 1496 1556 1504
rect 3372 1496 3380 1504
rect 3436 1496 3444 1504
rect 3628 1496 3636 1504
rect 3724 1496 3732 1504
rect 5548 1496 5556 1504
rect 7244 1496 7252 1504
rect 1100 1476 1108 1484
rect 2412 1476 2420 1484
rect 4300 1476 4308 1484
rect 4588 1476 4596 1484
rect 4652 1476 4660 1484
rect 4748 1476 4756 1484
rect 4876 1476 4884 1484
rect 5292 1476 5300 1484
rect 44 1456 52 1464
rect 1260 1456 1268 1464
rect 2764 1456 2772 1464
rect 4940 1456 4948 1464
rect 108 1436 116 1444
rect 1580 1436 1588 1444
rect 1676 1436 1684 1444
rect 1708 1436 1716 1444
rect 2540 1436 2548 1444
rect 3180 1436 3188 1444
rect 4076 1436 4084 1444
rect 5260 1456 5268 1464
rect 7116 1476 7124 1484
rect 5612 1456 5620 1464
rect 6284 1456 6292 1464
rect 6444 1456 6452 1464
rect 6924 1436 6932 1444
rect 4300 1416 4308 1424
rect 4972 1416 4980 1424
rect 5644 1416 5652 1424
rect 6476 1416 6484 1424
rect 7148 1416 7156 1424
rect 2916 1406 2923 1414
rect 2923 1406 2924 1414
rect 2928 1406 2933 1414
rect 2933 1406 2935 1414
rect 2935 1406 2936 1414
rect 2940 1406 2943 1414
rect 2943 1406 2945 1414
rect 2945 1406 2948 1414
rect 2952 1406 2953 1414
rect 2953 1406 2955 1414
rect 2955 1406 2960 1414
rect 2964 1406 2965 1414
rect 2965 1406 2972 1414
rect 5924 1406 5931 1414
rect 5931 1406 5932 1414
rect 5936 1406 5941 1414
rect 5941 1406 5943 1414
rect 5943 1406 5944 1414
rect 5948 1406 5951 1414
rect 5951 1406 5953 1414
rect 5953 1406 5956 1414
rect 5960 1406 5961 1414
rect 5961 1406 5963 1414
rect 5963 1406 5968 1414
rect 5972 1406 5973 1414
rect 5973 1406 5980 1414
rect 1228 1396 1236 1404
rect 1260 1396 1268 1404
rect 3084 1396 3092 1404
rect 3628 1396 3636 1404
rect 3820 1396 3828 1404
rect 5452 1396 5460 1404
rect 396 1376 404 1384
rect 1004 1356 1012 1364
rect 4236 1376 4244 1384
rect 4684 1376 4692 1384
rect 5548 1376 5556 1384
rect 6476 1376 6484 1384
rect 4940 1356 4948 1364
rect 6604 1356 6612 1364
rect 140 1336 148 1344
rect 2508 1336 2516 1344
rect 2604 1336 2612 1344
rect 3052 1336 3060 1344
rect 3340 1336 3348 1344
rect 3788 1336 3796 1344
rect 780 1316 788 1324
rect 2412 1316 2420 1324
rect 6220 1336 6228 1344
rect 6828 1336 6836 1344
rect 6924 1336 6932 1344
rect 4556 1316 4564 1324
rect 6796 1316 6804 1324
rect 6892 1316 6900 1324
rect 1004 1296 1012 1304
rect 1548 1296 1556 1304
rect 2508 1296 2516 1304
rect 4652 1296 4660 1304
rect 5292 1296 5300 1304
rect 6252 1296 6260 1304
rect 6604 1296 6612 1304
rect 3244 1276 3252 1284
rect 5100 1276 5108 1284
rect 6092 1276 6100 1284
rect 972 1256 980 1264
rect 1004 1256 1012 1264
rect 2348 1256 2356 1264
rect 3212 1256 3220 1264
rect 3436 1256 3444 1264
rect 5196 1256 5204 1264
rect 6028 1256 6036 1264
rect 1324 1236 1332 1244
rect 3596 1236 3604 1244
rect 4556 1236 4564 1244
rect 6188 1236 6196 1244
rect 1708 1216 1716 1224
rect 1900 1216 1908 1224
rect 3948 1216 3956 1224
rect 1412 1206 1419 1214
rect 1419 1206 1420 1214
rect 1424 1206 1429 1214
rect 1429 1206 1431 1214
rect 1431 1206 1432 1214
rect 1436 1206 1439 1214
rect 1439 1206 1441 1214
rect 1441 1206 1444 1214
rect 1448 1206 1449 1214
rect 1449 1206 1451 1214
rect 1451 1206 1456 1214
rect 1460 1206 1461 1214
rect 1461 1206 1468 1214
rect 4420 1206 4427 1214
rect 4427 1206 4428 1214
rect 4432 1206 4437 1214
rect 4437 1206 4439 1214
rect 4439 1206 4440 1214
rect 4444 1206 4447 1214
rect 4447 1206 4449 1214
rect 4449 1206 4452 1214
rect 4456 1206 4457 1214
rect 4457 1206 4459 1214
rect 4459 1206 4464 1214
rect 4468 1206 4469 1214
rect 4469 1206 4476 1214
rect 1580 1196 1588 1204
rect 2476 1196 2484 1204
rect 3500 1196 3508 1204
rect 1004 1176 1012 1184
rect 1676 1156 1684 1164
rect 364 1136 372 1144
rect 3948 1156 3956 1164
rect 4172 1156 4180 1164
rect 1036 1116 1044 1124
rect 236 1096 244 1104
rect 396 1096 404 1104
rect 2860 1116 2868 1124
rect 3468 1116 3476 1124
rect 4108 1116 4116 1124
rect 4364 1116 4372 1124
rect 5196 1136 5204 1144
rect 5452 1136 5460 1144
rect 6284 1136 6292 1144
rect 4908 1116 4916 1124
rect 5132 1116 5140 1124
rect 6476 1116 6484 1124
rect 6956 1116 6964 1124
rect 7052 1116 7060 1124
rect 2316 1096 2324 1104
rect 4204 1096 4212 1104
rect 4524 1096 4532 1104
rect 1036 1076 1044 1084
rect 1356 1076 1364 1084
rect 1676 1056 1684 1064
rect 2124 1056 2132 1064
rect 2540 1056 2548 1064
rect 3532 1076 3540 1084
rect 4172 1076 4180 1084
rect 5068 1096 5076 1104
rect 5324 1096 5332 1104
rect 4620 1076 4628 1084
rect 6188 1096 6196 1104
rect 5612 1076 5620 1084
rect 7308 1076 7316 1084
rect 108 1036 116 1044
rect 4076 1056 4084 1064
rect 4524 1056 4532 1064
rect 6188 1036 6196 1044
rect 7308 1036 7316 1044
rect 3020 1016 3028 1024
rect 4044 1016 4052 1024
rect 6028 1016 6036 1024
rect 7372 1016 7380 1024
rect 2916 1006 2923 1014
rect 2923 1006 2924 1014
rect 2928 1006 2933 1014
rect 2933 1006 2935 1014
rect 2935 1006 2936 1014
rect 2940 1006 2943 1014
rect 2943 1006 2945 1014
rect 2945 1006 2948 1014
rect 2952 1006 2953 1014
rect 2953 1006 2955 1014
rect 2955 1006 2960 1014
rect 2964 1006 2965 1014
rect 2965 1006 2972 1014
rect 5924 1006 5931 1014
rect 5931 1006 5932 1014
rect 5936 1006 5941 1014
rect 5941 1006 5943 1014
rect 5943 1006 5944 1014
rect 5948 1006 5951 1014
rect 5951 1006 5953 1014
rect 5953 1006 5956 1014
rect 5960 1006 5961 1014
rect 5961 1006 5963 1014
rect 5963 1006 5968 1014
rect 5972 1006 5973 1014
rect 5973 1006 5980 1014
rect 748 996 756 1004
rect 1100 996 1108 1004
rect 2092 976 2100 984
rect 2220 976 2228 984
rect 3660 996 3668 1004
rect 3372 976 3380 984
rect 7308 996 7316 1004
rect 7372 976 7380 984
rect 1292 936 1300 944
rect 3116 956 3124 964
rect 3372 936 3380 944
rect 7116 956 7124 964
rect 5452 936 5460 944
rect 236 916 244 924
rect 2060 916 2068 924
rect 2092 916 2100 924
rect 2220 916 2228 924
rect 4780 916 4788 924
rect 5772 916 5780 924
rect 7244 916 7252 924
rect 4748 896 4756 904
rect 1292 876 1300 884
rect 1612 876 1620 884
rect 1900 876 1908 884
rect 2060 876 2068 884
rect 2124 876 2132 884
rect 4588 876 4596 884
rect 5804 896 5812 904
rect 6252 896 6260 904
rect 7276 896 7284 904
rect 780 856 788 864
rect 2572 856 2580 864
rect 1260 836 1268 844
rect 6444 856 6452 864
rect 6668 836 6676 844
rect 3980 816 3988 824
rect 1412 806 1419 814
rect 1419 806 1420 814
rect 1424 806 1429 814
rect 1429 806 1431 814
rect 1431 806 1432 814
rect 1436 806 1439 814
rect 1439 806 1441 814
rect 1441 806 1444 814
rect 1448 806 1449 814
rect 1449 806 1451 814
rect 1451 806 1456 814
rect 1460 806 1461 814
rect 1461 806 1468 814
rect 4420 806 4427 814
rect 4427 806 4428 814
rect 4432 806 4437 814
rect 4437 806 4439 814
rect 4439 806 4440 814
rect 4444 806 4447 814
rect 4447 806 4449 814
rect 4449 806 4452 814
rect 4456 806 4457 814
rect 4457 806 4459 814
rect 4459 806 4464 814
rect 4468 806 4469 814
rect 4469 806 4476 814
rect 4844 796 4852 804
rect 1868 776 1876 784
rect 4236 776 4244 784
rect 4876 776 4884 784
rect 6700 776 6708 784
rect 844 756 852 764
rect 1036 756 1044 764
rect 2444 756 2452 764
rect 4044 756 4052 764
rect 2316 736 2324 744
rect 1164 716 1172 724
rect 4332 736 4340 744
rect 6284 736 6292 744
rect 7084 736 7092 744
rect 2860 716 2868 724
rect 3948 716 3956 724
rect 4940 716 4948 724
rect 5804 716 5812 724
rect 2284 696 2292 704
rect 3852 696 3860 704
rect 6028 696 6036 704
rect 6284 696 6292 704
rect 6700 696 6708 704
rect 140 676 148 684
rect 1004 676 1012 684
rect 2156 676 2164 684
rect 4236 676 4244 684
rect 4780 676 4788 684
rect 4876 676 4884 684
rect 7212 676 7220 684
rect 2284 656 2292 664
rect 2540 656 2548 664
rect 4044 656 4052 664
rect 5036 656 5044 664
rect 7340 656 7348 664
rect 812 636 820 644
rect 3756 636 3764 644
rect 4204 636 4212 644
rect 2476 616 2484 624
rect 2916 606 2923 614
rect 2923 606 2924 614
rect 2928 606 2933 614
rect 2933 606 2935 614
rect 2935 606 2936 614
rect 2940 606 2943 614
rect 2943 606 2945 614
rect 2945 606 2948 614
rect 2952 606 2953 614
rect 2953 606 2955 614
rect 2955 606 2960 614
rect 2964 606 2965 614
rect 2965 606 2972 614
rect 4108 616 4116 624
rect 4972 616 4980 624
rect 5772 616 5780 624
rect 6604 636 6612 644
rect 7308 636 7316 644
rect 5924 606 5931 614
rect 5931 606 5932 614
rect 5936 606 5941 614
rect 5941 606 5943 614
rect 5943 606 5944 614
rect 5948 606 5951 614
rect 5951 606 5953 614
rect 5953 606 5956 614
rect 5960 606 5961 614
rect 5961 606 5963 614
rect 5963 606 5968 614
rect 5972 606 5973 614
rect 5973 606 5980 614
rect 5196 596 5204 604
rect 5612 596 5620 604
rect 2476 576 2484 584
rect 4524 576 4532 584
rect 4812 576 4820 584
rect 6124 576 6132 584
rect 1164 556 1172 564
rect 748 536 756 544
rect 2156 536 2164 544
rect 3596 536 3604 544
rect 3948 536 3956 544
rect 3980 536 3988 544
rect 4652 536 4660 544
rect 5004 536 5012 544
rect 7116 536 7124 544
rect 1868 516 1876 524
rect 4364 516 4372 524
rect 4748 516 4756 524
rect 4908 516 4916 524
rect 5804 516 5812 524
rect 44 496 52 504
rect 140 496 148 504
rect 1324 496 1332 504
rect 1740 496 1748 504
rect 2188 496 2196 504
rect 6476 496 6484 504
rect 2444 476 2452 484
rect 2572 476 2580 484
rect 4172 476 4180 484
rect 6060 476 6068 484
rect 5804 456 5812 464
rect 7180 436 7188 444
rect 1412 406 1419 414
rect 1419 406 1420 414
rect 1424 406 1429 414
rect 1429 406 1431 414
rect 1431 406 1432 414
rect 1436 406 1439 414
rect 1439 406 1441 414
rect 1441 406 1444 414
rect 1448 406 1449 414
rect 1449 406 1451 414
rect 1451 406 1456 414
rect 1460 406 1461 414
rect 1461 406 1468 414
rect 4420 406 4427 414
rect 4427 406 4428 414
rect 4432 406 4437 414
rect 4437 406 4439 414
rect 4439 406 4440 414
rect 4444 406 4447 414
rect 4447 406 4449 414
rect 4449 406 4452 414
rect 4456 406 4457 414
rect 4457 406 4459 414
rect 4459 406 4464 414
rect 4468 406 4469 414
rect 4469 406 4476 414
rect 364 376 372 384
rect 3852 376 3860 384
rect 4300 356 4308 364
rect 1868 336 1876 344
rect 1964 336 1972 344
rect 3884 336 3892 344
rect 2092 316 2100 324
rect 2284 316 2292 324
rect 3212 316 3220 324
rect 6188 316 6196 324
rect 7404 316 7412 324
rect 780 296 788 304
rect 1164 296 1172 304
rect 844 276 852 284
rect 1836 276 1844 284
rect 1964 276 1972 284
rect 876 256 884 264
rect 4076 296 4084 304
rect 4812 296 4820 304
rect 4844 296 4852 304
rect 6796 296 6804 304
rect 7372 296 7380 304
rect 4044 276 4052 284
rect 4300 276 4308 284
rect 4620 276 4628 284
rect 5100 276 5108 284
rect 2092 256 2100 264
rect 3340 256 3348 264
rect 3180 236 3188 244
rect 4940 236 4948 244
rect 2916 206 2923 214
rect 2923 206 2924 214
rect 2928 206 2933 214
rect 2933 206 2935 214
rect 2935 206 2936 214
rect 2940 206 2943 214
rect 2943 206 2945 214
rect 2945 206 2948 214
rect 2952 206 2953 214
rect 2953 206 2955 214
rect 2955 206 2960 214
rect 2964 206 2965 214
rect 2965 206 2972 214
rect 5924 206 5931 214
rect 5931 206 5932 214
rect 5936 206 5941 214
rect 5941 206 5943 214
rect 5943 206 5944 214
rect 5948 206 5951 214
rect 5951 206 5953 214
rect 5953 206 5956 214
rect 5960 206 5961 214
rect 5961 206 5963 214
rect 5963 206 5968 214
rect 5972 206 5973 214
rect 5973 206 5980 214
rect 364 156 372 164
rect 1036 176 1044 184
rect 2284 176 2292 184
rect 3884 176 3892 184
rect 4620 176 4628 184
rect 4844 196 4852 204
rect 6668 176 6676 184
rect 6732 176 6740 184
rect 6924 176 6932 184
rect 812 156 820 164
rect 5036 156 5044 164
rect 6380 156 6388 164
rect 4652 136 4660 144
rect 7020 136 7028 144
rect 3756 96 3764 104
rect 4844 96 4852 104
rect 5068 96 5076 104
rect 6636 96 6644 104
rect 4876 76 4884 84
rect 4812 36 4820 44
rect 3468 16 3476 24
rect 3596 16 3604 24
rect 3660 16 3668 24
rect 4076 16 4084 24
rect 5196 16 5204 24
rect 1412 6 1419 14
rect 1419 6 1420 14
rect 1424 6 1429 14
rect 1429 6 1431 14
rect 1431 6 1432 14
rect 1436 6 1439 14
rect 1439 6 1441 14
rect 1441 6 1444 14
rect 1448 6 1449 14
rect 1449 6 1451 14
rect 1451 6 1456 14
rect 1460 6 1461 14
rect 1461 6 1468 14
rect 4420 6 4427 14
rect 4427 6 4428 14
rect 4432 6 4437 14
rect 4437 6 4439 14
rect 4439 6 4440 14
rect 4444 6 4447 14
rect 4447 6 4449 14
rect 4449 6 4452 14
rect 4456 6 4457 14
rect 4457 6 4459 14
rect 4459 6 4464 14
rect 4468 6 4469 14
rect 4469 6 4476 14
<< metal4 >>
rect 3434 5424 3446 5426
rect 3434 5416 3436 5424
rect 3444 5416 3446 5424
rect 1408 5214 1472 5416
rect 2912 5414 2976 5416
rect 2912 5406 2916 5414
rect 2924 5406 2928 5414
rect 2936 5406 2940 5414
rect 2948 5406 2952 5414
rect 2960 5406 2964 5414
rect 2972 5406 2976 5414
rect 1610 5344 1622 5346
rect 1610 5336 1612 5344
rect 1620 5336 1622 5344
rect 1610 5326 1622 5336
rect 1610 5314 1686 5326
rect 1674 5304 1686 5314
rect 1674 5296 1676 5304
rect 1684 5296 1686 5304
rect 1674 5294 1686 5296
rect 1408 5206 1412 5214
rect 1420 5206 1424 5214
rect 1432 5206 1436 5214
rect 1444 5206 1448 5214
rect 1456 5206 1460 5214
rect 1468 5206 1472 5214
rect 138 5144 150 5146
rect 138 5136 140 5144
rect 148 5136 150 5144
rect 106 4984 118 4986
rect 106 4976 108 4984
rect 116 4976 118 4984
rect 106 4284 118 4976
rect 138 4684 150 5136
rect 202 5104 214 5106
rect 202 5096 204 5104
rect 212 5096 214 5104
rect 202 4964 214 5096
rect 1322 5104 1334 5106
rect 1322 5096 1324 5104
rect 1332 5096 1334 5104
rect 970 5024 982 5026
rect 970 5016 972 5024
rect 980 5016 982 5024
rect 202 4956 204 4964
rect 212 4956 214 4964
rect 202 4954 214 4956
rect 330 4964 342 4966
rect 330 4956 332 4964
rect 340 4956 342 4964
rect 138 4676 140 4684
rect 148 4676 150 4684
rect 138 4674 150 4676
rect 298 4684 310 4686
rect 298 4676 300 4684
rect 308 4676 310 4684
rect 106 4276 108 4284
rect 116 4276 118 4284
rect 106 4274 118 4276
rect 10 3964 22 3966
rect 10 3956 12 3964
rect 20 3956 22 3964
rect 10 3764 22 3956
rect 10 3756 12 3764
rect 20 3756 22 3764
rect 10 3754 22 3756
rect 170 3924 182 3926
rect 170 3916 172 3924
rect 180 3916 182 3924
rect 170 3724 182 3916
rect 170 3716 172 3724
rect 180 3716 182 3724
rect 170 3714 182 3716
rect 298 3544 310 4676
rect 298 3536 300 3544
rect 308 3536 310 3544
rect 298 3534 310 3536
rect 330 3484 342 4956
rect 970 4844 982 5016
rect 1258 4964 1286 4966
rect 1258 4956 1276 4964
rect 1284 4956 1286 4964
rect 1258 4954 1286 4956
rect 1258 4924 1270 4954
rect 1258 4916 1260 4924
rect 1268 4916 1270 4924
rect 1258 4914 1270 4916
rect 1322 4904 1334 5096
rect 1322 4896 1324 4904
rect 1332 4896 1334 4904
rect 1322 4894 1334 4896
rect 970 4836 972 4844
rect 980 4836 982 4844
rect 970 4834 982 4836
rect 1354 4864 1366 4866
rect 1354 4856 1356 4864
rect 1364 4856 1366 4864
rect 1322 4744 1334 4746
rect 1322 4736 1324 4744
rect 1332 4736 1334 4744
rect 842 4724 854 4726
rect 842 4716 844 4724
rect 852 4716 854 4724
rect 778 4384 790 4386
rect 778 4376 780 4384
rect 788 4376 790 4384
rect 746 4364 758 4366
rect 746 4356 748 4364
rect 756 4356 758 4364
rect 522 4324 534 4326
rect 522 4316 524 4324
rect 532 4316 534 4324
rect 330 3476 332 3484
rect 340 3476 342 3484
rect 330 3474 342 3476
rect 394 3944 406 3946
rect 394 3936 396 3944
rect 404 3936 406 3944
rect 202 3124 214 3126
rect 202 3116 204 3124
rect 212 3116 214 3124
rect 74 3104 86 3106
rect 74 3096 76 3104
rect 84 3096 86 3104
rect 74 1724 86 3096
rect 170 2364 182 2366
rect 170 2356 172 2364
rect 180 2356 182 2364
rect 170 2064 182 2356
rect 170 2056 172 2064
rect 180 2056 182 2064
rect 170 2054 182 2056
rect 74 1716 76 1724
rect 84 1716 86 1724
rect 74 1714 86 1716
rect 138 1844 150 1846
rect 138 1836 140 1844
rect 148 1836 150 1844
rect 42 1464 54 1466
rect 42 1456 44 1464
rect 52 1456 54 1464
rect 42 504 54 1456
rect 106 1444 118 1446
rect 106 1436 108 1444
rect 116 1436 118 1444
rect 106 1044 118 1436
rect 138 1344 150 1836
rect 202 1724 214 3116
rect 394 3124 406 3936
rect 522 3664 534 4316
rect 522 3656 524 3664
rect 532 3656 534 3664
rect 522 3654 534 3656
rect 650 3724 662 3726
rect 650 3716 652 3724
rect 660 3716 662 3724
rect 650 3324 662 3716
rect 746 3524 758 4356
rect 778 4144 790 4376
rect 778 4136 780 4144
rect 788 4136 790 4144
rect 778 4134 790 4136
rect 810 3804 822 3806
rect 810 3796 812 3804
rect 820 3796 822 3804
rect 810 3724 822 3796
rect 810 3716 812 3724
rect 820 3716 822 3724
rect 810 3714 822 3716
rect 842 3644 854 4716
rect 1290 4584 1302 4586
rect 1290 4576 1292 4584
rect 1300 4576 1302 4584
rect 874 4324 886 4326
rect 874 4316 876 4324
rect 884 4316 886 4324
rect 874 3764 886 4316
rect 1226 4324 1238 4326
rect 1226 4316 1228 4324
rect 1236 4316 1238 4324
rect 1066 4304 1078 4306
rect 1066 4296 1068 4304
rect 1076 4296 1078 4304
rect 906 4284 918 4286
rect 906 4276 908 4284
rect 916 4276 918 4284
rect 906 3904 918 4276
rect 1002 4244 1014 4246
rect 1002 4236 1004 4244
rect 1012 4236 1014 4244
rect 906 3896 908 3904
rect 916 3896 918 3904
rect 906 3894 918 3896
rect 970 4204 982 4206
rect 970 4196 972 4204
rect 980 4196 982 4204
rect 874 3756 876 3764
rect 884 3756 886 3764
rect 874 3754 886 3756
rect 970 3864 982 4196
rect 970 3856 972 3864
rect 980 3856 982 3864
rect 842 3636 844 3644
rect 852 3636 854 3644
rect 842 3634 854 3636
rect 906 3724 918 3726
rect 906 3716 908 3724
rect 916 3716 918 3724
rect 746 3516 748 3524
rect 756 3516 758 3524
rect 746 3514 758 3516
rect 650 3316 652 3324
rect 660 3316 662 3324
rect 650 3314 662 3316
rect 714 3504 726 3506
rect 714 3496 716 3504
rect 724 3496 726 3504
rect 394 3116 396 3124
rect 404 3116 406 3124
rect 394 3114 406 3116
rect 714 3124 726 3496
rect 874 3504 886 3506
rect 874 3496 876 3504
rect 884 3496 886 3504
rect 874 3404 886 3496
rect 874 3396 876 3404
rect 884 3396 886 3404
rect 778 3364 790 3366
rect 778 3356 780 3364
rect 788 3356 790 3364
rect 714 3116 716 3124
rect 724 3116 726 3124
rect 714 3114 726 3116
rect 746 3124 758 3126
rect 746 3116 748 3124
rect 756 3116 758 3124
rect 362 3104 374 3106
rect 362 3096 364 3104
rect 372 3096 374 3104
rect 362 2864 374 3096
rect 362 2856 364 2864
rect 372 2856 374 2864
rect 362 2854 374 2856
rect 554 3104 566 3106
rect 554 3096 556 3104
rect 564 3096 566 3104
rect 554 2704 566 3096
rect 586 3084 598 3086
rect 586 3076 588 3084
rect 596 3076 598 3084
rect 586 2904 598 3076
rect 586 2896 588 2904
rect 596 2896 598 2904
rect 586 2894 598 2896
rect 714 3084 726 3086
rect 714 3076 716 3084
rect 724 3076 726 3084
rect 554 2696 556 2704
rect 564 2696 566 2704
rect 554 2694 566 2696
rect 650 2744 662 2746
rect 650 2736 652 2744
rect 660 2736 662 2744
rect 362 2684 374 2686
rect 362 2676 364 2684
rect 372 2676 374 2684
rect 202 1716 204 1724
rect 212 1716 214 1724
rect 202 1714 214 1716
rect 266 1764 278 1766
rect 266 1756 268 1764
rect 276 1756 278 1764
rect 266 1724 278 1756
rect 266 1716 268 1724
rect 276 1716 278 1724
rect 266 1714 278 1716
rect 138 1336 140 1344
rect 148 1336 150 1344
rect 138 1334 150 1336
rect 362 1144 374 2676
rect 458 2564 470 2566
rect 458 2556 460 2564
rect 468 2556 470 2564
rect 458 2284 470 2556
rect 458 2276 460 2284
rect 468 2276 470 2284
rect 458 2274 470 2276
rect 522 2124 534 2126
rect 522 2116 524 2124
rect 532 2116 534 2124
rect 522 1884 534 2116
rect 650 2124 662 2736
rect 650 2116 652 2124
rect 660 2116 662 2124
rect 650 2114 662 2116
rect 682 2304 694 2306
rect 682 2296 684 2304
rect 692 2296 694 2304
rect 522 1876 524 1884
rect 532 1876 534 1884
rect 522 1874 534 1876
rect 682 1744 694 2296
rect 714 2044 726 3076
rect 746 2744 758 3116
rect 778 3084 790 3356
rect 778 3076 780 3084
rect 788 3076 790 3084
rect 778 3074 790 3076
rect 810 3004 822 3006
rect 810 2996 812 3004
rect 820 2996 822 3004
rect 746 2736 748 2744
rect 756 2736 758 2744
rect 746 2734 758 2736
rect 778 2784 790 2786
rect 778 2776 780 2784
rect 788 2776 790 2784
rect 778 2484 790 2776
rect 810 2644 822 2996
rect 874 2784 886 3396
rect 906 3024 918 3716
rect 970 3684 982 3856
rect 970 3676 972 3684
rect 980 3676 982 3684
rect 970 3674 982 3676
rect 1002 3844 1014 4236
rect 1034 4184 1046 4186
rect 1034 4176 1036 4184
rect 1044 4176 1046 4184
rect 1034 3924 1046 4176
rect 1066 4104 1078 4296
rect 1066 4096 1068 4104
rect 1076 4096 1078 4104
rect 1066 4094 1078 4096
rect 1162 4144 1174 4146
rect 1162 4136 1164 4144
rect 1172 4136 1174 4144
rect 1162 4104 1174 4136
rect 1162 4096 1164 4104
rect 1172 4096 1174 4104
rect 1162 4094 1174 4096
rect 1034 3916 1036 3924
rect 1044 3916 1046 3924
rect 1034 3914 1046 3916
rect 1002 3836 1004 3844
rect 1012 3836 1014 3844
rect 906 3016 908 3024
rect 916 3016 918 3024
rect 906 3014 918 3016
rect 874 2776 876 2784
rect 884 2776 886 2784
rect 874 2774 886 2776
rect 810 2636 812 2644
rect 820 2636 822 2644
rect 810 2634 822 2636
rect 842 2644 854 2646
rect 842 2636 844 2644
rect 852 2636 854 2644
rect 778 2476 780 2484
rect 788 2476 790 2484
rect 778 2474 790 2476
rect 714 2036 716 2044
rect 724 2036 726 2044
rect 714 2034 726 2036
rect 778 2344 790 2346
rect 778 2336 780 2344
rect 788 2336 790 2344
rect 778 1964 790 2336
rect 778 1956 780 1964
rect 788 1956 790 1964
rect 778 1954 790 1956
rect 682 1736 684 1744
rect 692 1736 694 1744
rect 682 1734 694 1736
rect 362 1136 364 1144
rect 372 1136 374 1144
rect 362 1134 374 1136
rect 394 1384 406 1386
rect 394 1376 396 1384
rect 404 1376 406 1384
rect 106 1036 108 1044
rect 116 1036 118 1044
rect 106 1034 118 1036
rect 234 1104 246 1106
rect 234 1096 236 1104
rect 244 1096 246 1104
rect 234 924 246 1096
rect 394 1104 406 1376
rect 394 1096 396 1104
rect 404 1096 406 1104
rect 394 1094 406 1096
rect 778 1324 790 1326
rect 778 1316 780 1324
rect 788 1316 790 1324
rect 234 916 236 924
rect 244 916 246 924
rect 234 914 246 916
rect 746 1004 758 1006
rect 746 996 748 1004
rect 756 996 758 1004
rect 42 496 44 504
rect 52 496 54 504
rect 42 494 54 496
rect 138 684 150 686
rect 138 676 140 684
rect 148 676 150 684
rect 138 504 150 676
rect 746 544 758 996
rect 746 536 748 544
rect 756 536 758 544
rect 746 534 758 536
rect 778 864 790 1316
rect 778 856 780 864
rect 788 856 790 864
rect 138 496 140 504
rect 148 496 150 504
rect 138 494 150 496
rect 362 384 374 386
rect 362 376 364 384
rect 372 376 374 384
rect 362 164 374 376
rect 778 304 790 856
rect 842 764 854 2636
rect 1002 2424 1014 3836
rect 1034 3784 1046 3786
rect 1034 3776 1036 3784
rect 1044 3776 1046 3784
rect 1034 3324 1046 3776
rect 1226 3544 1238 4316
rect 1290 3924 1302 4576
rect 1322 4064 1334 4736
rect 1322 4056 1324 4064
rect 1332 4056 1334 4064
rect 1322 4054 1334 4056
rect 1354 3984 1366 4856
rect 1354 3976 1356 3984
rect 1364 3976 1366 3984
rect 1354 3974 1366 3976
rect 1408 4814 1472 5206
rect 1898 5184 1910 5186
rect 1898 5176 1900 5184
rect 1908 5176 1910 5184
rect 1770 5104 1782 5106
rect 1770 5096 1772 5104
rect 1780 5096 1782 5104
rect 1408 4806 1412 4814
rect 1420 4806 1424 4814
rect 1432 4806 1436 4814
rect 1444 4806 1448 4814
rect 1456 4806 1460 4814
rect 1468 4806 1472 4814
rect 1408 4414 1472 4806
rect 1578 4964 1590 4966
rect 1578 4956 1580 4964
rect 1588 4956 1590 4964
rect 1578 4484 1590 4956
rect 1770 4924 1782 5096
rect 1898 4964 1910 5176
rect 2666 5184 2678 5186
rect 2666 5176 2668 5184
rect 2676 5176 2678 5184
rect 2570 5024 2582 5026
rect 2570 5016 2572 5024
rect 2580 5016 2582 5024
rect 1898 4956 1900 4964
rect 1908 4956 1910 4964
rect 1898 4954 1910 4956
rect 2026 4984 2038 4986
rect 2026 4976 2028 4984
rect 2036 4976 2038 4984
rect 1770 4916 1772 4924
rect 1780 4916 1782 4924
rect 1770 4914 1782 4916
rect 2026 4864 2038 4976
rect 2410 4984 2422 4986
rect 2410 4976 2412 4984
rect 2420 4976 2422 4984
rect 2250 4944 2262 4946
rect 2250 4936 2252 4944
rect 2260 4936 2262 4944
rect 2026 4856 2028 4864
rect 2036 4856 2038 4864
rect 2026 4854 2038 4856
rect 2058 4924 2070 4926
rect 2058 4916 2060 4924
rect 2068 4916 2070 4924
rect 2058 4864 2070 4916
rect 2058 4856 2060 4864
rect 2068 4856 2070 4864
rect 2058 4854 2070 4856
rect 1674 4764 1686 4766
rect 1674 4756 1676 4764
rect 1684 4756 1686 4764
rect 1578 4476 1580 4484
rect 1588 4476 1590 4484
rect 1578 4474 1590 4476
rect 1642 4704 1654 4706
rect 1642 4696 1644 4704
rect 1652 4696 1654 4704
rect 1642 4464 1654 4696
rect 1642 4456 1644 4464
rect 1652 4456 1654 4464
rect 1642 4454 1654 4456
rect 1408 4406 1412 4414
rect 1420 4406 1424 4414
rect 1432 4406 1436 4414
rect 1444 4406 1448 4414
rect 1456 4406 1460 4414
rect 1468 4406 1472 4414
rect 1408 4014 1472 4406
rect 1578 4304 1590 4306
rect 1578 4296 1580 4304
rect 1588 4296 1590 4304
rect 1408 4006 1412 4014
rect 1420 4006 1424 4014
rect 1432 4006 1436 4014
rect 1444 4006 1448 4014
rect 1456 4006 1460 4014
rect 1468 4006 1472 4014
rect 1290 3916 1292 3924
rect 1300 3916 1302 3924
rect 1290 3914 1302 3916
rect 1354 3944 1366 3946
rect 1354 3936 1356 3944
rect 1364 3936 1366 3944
rect 1226 3536 1228 3544
rect 1236 3536 1238 3544
rect 1226 3534 1238 3536
rect 1290 3804 1302 3806
rect 1290 3796 1292 3804
rect 1300 3796 1302 3804
rect 1034 3316 1036 3324
rect 1044 3316 1046 3324
rect 1034 3314 1046 3316
rect 1034 3064 1046 3066
rect 1034 3056 1036 3064
rect 1044 3056 1046 3064
rect 1034 2924 1046 3056
rect 1034 2916 1036 2924
rect 1044 2916 1046 2924
rect 1034 2914 1046 2916
rect 1290 2924 1302 3796
rect 1354 3744 1366 3936
rect 1354 3736 1356 3744
rect 1364 3736 1366 3744
rect 1354 3734 1366 3736
rect 1408 3614 1472 4006
rect 1408 3606 1412 3614
rect 1420 3606 1424 3614
rect 1432 3606 1436 3614
rect 1444 3606 1448 3614
rect 1456 3606 1460 3614
rect 1468 3606 1472 3614
rect 1290 2916 1292 2924
rect 1300 2916 1302 2924
rect 1290 2914 1302 2916
rect 1354 3344 1366 3346
rect 1354 3336 1356 3344
rect 1364 3336 1366 3344
rect 1354 2884 1366 3336
rect 1354 2876 1356 2884
rect 1364 2876 1366 2884
rect 1354 2874 1366 2876
rect 1408 3214 1472 3606
rect 1408 3206 1412 3214
rect 1420 3206 1424 3214
rect 1432 3206 1436 3214
rect 1444 3206 1448 3214
rect 1456 3206 1460 3214
rect 1468 3206 1472 3214
rect 1408 2814 1472 3206
rect 1514 4064 1526 4066
rect 1514 4056 1516 4064
rect 1524 4056 1526 4064
rect 1514 3164 1526 4056
rect 1546 3904 1558 3906
rect 1546 3896 1548 3904
rect 1556 3896 1558 3904
rect 1546 3184 1558 3896
rect 1546 3176 1548 3184
rect 1556 3176 1558 3184
rect 1546 3174 1558 3176
rect 1514 3156 1516 3164
rect 1524 3156 1526 3164
rect 1514 3154 1526 3156
rect 1408 2806 1412 2814
rect 1420 2806 1424 2814
rect 1432 2806 1436 2814
rect 1444 2806 1448 2814
rect 1456 2806 1460 2814
rect 1468 2806 1472 2814
rect 1130 2704 1142 2706
rect 1130 2696 1132 2704
rect 1140 2696 1142 2704
rect 1002 2416 1004 2424
rect 1012 2416 1014 2424
rect 1002 2414 1014 2416
rect 1098 2424 1110 2426
rect 1098 2416 1100 2424
rect 1108 2416 1110 2424
rect 970 2344 982 2346
rect 970 2336 972 2344
rect 980 2336 982 2344
rect 938 1784 950 1786
rect 938 1776 940 1784
rect 948 1776 950 1784
rect 938 1504 950 1776
rect 970 1744 982 2336
rect 970 1736 972 1744
rect 980 1736 982 1744
rect 970 1684 982 1736
rect 1002 1844 1014 1846
rect 1002 1836 1004 1844
rect 1012 1836 1014 1844
rect 1002 1724 1014 1836
rect 1002 1716 1004 1724
rect 1012 1716 1014 1724
rect 1002 1714 1014 1716
rect 970 1676 972 1684
rect 980 1676 982 1684
rect 970 1674 982 1676
rect 938 1496 940 1504
rect 948 1496 950 1504
rect 938 1494 950 1496
rect 970 1544 982 1546
rect 970 1536 972 1544
rect 980 1536 982 1544
rect 970 1264 982 1536
rect 1098 1524 1110 2416
rect 1130 2224 1142 2696
rect 1162 2704 1174 2706
rect 1162 2696 1164 2704
rect 1172 2696 1174 2704
rect 1162 2264 1174 2696
rect 1258 2704 1270 2706
rect 1258 2696 1260 2704
rect 1268 2696 1270 2704
rect 1162 2256 1164 2264
rect 1172 2256 1174 2264
rect 1162 2254 1174 2256
rect 1226 2664 1238 2666
rect 1226 2656 1228 2664
rect 1236 2656 1238 2664
rect 1130 2216 1132 2224
rect 1140 2216 1142 2224
rect 1130 1804 1142 2216
rect 1194 2204 1206 2206
rect 1194 2196 1196 2204
rect 1204 2196 1206 2204
rect 1194 2004 1206 2196
rect 1226 2104 1238 2656
rect 1258 2304 1270 2696
rect 1322 2504 1334 2506
rect 1322 2496 1324 2504
rect 1332 2496 1334 2504
rect 1322 2424 1334 2496
rect 1322 2416 1324 2424
rect 1332 2416 1334 2424
rect 1322 2414 1334 2416
rect 1408 2414 1472 2806
rect 1408 2406 1412 2414
rect 1420 2406 1424 2414
rect 1432 2406 1436 2414
rect 1444 2406 1448 2414
rect 1456 2406 1460 2414
rect 1468 2406 1472 2414
rect 1258 2296 1260 2304
rect 1268 2296 1270 2304
rect 1258 2294 1270 2296
rect 1354 2304 1366 2306
rect 1354 2296 1356 2304
rect 1364 2296 1366 2304
rect 1226 2096 1228 2104
rect 1236 2096 1238 2104
rect 1226 2094 1238 2096
rect 1290 2284 1302 2286
rect 1290 2276 1292 2284
rect 1300 2276 1302 2284
rect 1258 2064 1270 2066
rect 1258 2056 1260 2064
rect 1268 2056 1270 2064
rect 1194 1996 1196 2004
rect 1204 1996 1206 2004
rect 1194 1994 1206 1996
rect 1226 2044 1238 2046
rect 1226 2036 1228 2044
rect 1236 2036 1238 2044
rect 1130 1796 1132 1804
rect 1140 1796 1142 1804
rect 1130 1724 1142 1796
rect 1130 1716 1132 1724
rect 1140 1716 1142 1724
rect 1130 1714 1142 1716
rect 1098 1516 1100 1524
rect 1108 1516 1110 1524
rect 1098 1514 1110 1516
rect 1098 1484 1110 1486
rect 1098 1476 1100 1484
rect 1108 1476 1110 1484
rect 1002 1364 1014 1366
rect 1002 1356 1004 1364
rect 1012 1356 1014 1364
rect 1002 1304 1014 1356
rect 1002 1296 1004 1304
rect 1012 1296 1014 1304
rect 1002 1294 1014 1296
rect 970 1256 972 1264
rect 980 1256 982 1264
rect 970 1254 982 1256
rect 1002 1264 1014 1266
rect 1002 1256 1004 1264
rect 1012 1256 1014 1264
rect 842 756 844 764
rect 852 756 854 764
rect 842 754 854 756
rect 1002 1184 1014 1256
rect 1002 1176 1004 1184
rect 1012 1176 1014 1184
rect 1002 684 1014 1176
rect 1034 1124 1046 1126
rect 1034 1116 1036 1124
rect 1044 1116 1046 1124
rect 1034 1084 1046 1116
rect 1034 1076 1036 1084
rect 1044 1076 1046 1084
rect 1034 1074 1046 1076
rect 1098 1004 1110 1476
rect 1226 1404 1238 2036
rect 1258 1464 1270 2056
rect 1290 1784 1302 2276
rect 1354 2164 1366 2296
rect 1354 2156 1356 2164
rect 1364 2156 1366 2164
rect 1354 2154 1366 2156
rect 1290 1776 1292 1784
rect 1300 1776 1302 1784
rect 1290 1774 1302 1776
rect 1322 2144 1334 2146
rect 1322 2136 1324 2144
rect 1332 2136 1334 2144
rect 1322 1764 1334 2136
rect 1408 2014 1472 2406
rect 1408 2006 1412 2014
rect 1420 2006 1424 2014
rect 1432 2006 1436 2014
rect 1444 2006 1448 2014
rect 1456 2006 1460 2014
rect 1468 2006 1472 2014
rect 1322 1756 1324 1764
rect 1332 1756 1334 1764
rect 1322 1754 1334 1756
rect 1354 1764 1366 1766
rect 1354 1756 1356 1764
rect 1364 1756 1366 1764
rect 1354 1684 1366 1756
rect 1354 1676 1356 1684
rect 1364 1676 1366 1684
rect 1354 1674 1366 1676
rect 1408 1614 1472 2006
rect 1514 2784 1526 2786
rect 1514 2776 1516 2784
rect 1524 2776 1526 2784
rect 1514 1624 1526 2776
rect 1578 2784 1590 4296
rect 1642 3984 1654 3986
rect 1642 3976 1644 3984
rect 1652 3976 1654 3984
rect 1642 3604 1654 3976
rect 1674 3944 1686 4756
rect 1962 4724 1974 4726
rect 1962 4716 1964 4724
rect 1972 4716 1974 4724
rect 1962 4604 1974 4716
rect 1962 4596 1964 4604
rect 1972 4596 1974 4604
rect 1962 4594 1974 4596
rect 1674 3936 1676 3944
rect 1684 3936 1686 3944
rect 1674 3934 1686 3936
rect 1706 4544 1718 4546
rect 1706 4536 1708 4544
rect 1716 4536 1718 4544
rect 1706 4284 1718 4536
rect 2122 4304 2134 4306
rect 2122 4296 2124 4304
rect 2132 4296 2134 4304
rect 1706 4276 1708 4284
rect 1716 4276 1718 4284
rect 1706 3924 1718 4276
rect 1770 4284 1782 4286
rect 1770 4276 1772 4284
rect 1780 4276 1782 4284
rect 1770 4244 1782 4276
rect 1770 4236 1772 4244
rect 1780 4236 1782 4244
rect 1770 4234 1782 4236
rect 1706 3916 1708 3924
rect 1716 3916 1718 3924
rect 1706 3914 1718 3916
rect 1642 3596 1644 3604
rect 1652 3596 1654 3604
rect 1642 3594 1654 3596
rect 1674 3904 1686 3906
rect 1674 3896 1676 3904
rect 1684 3896 1686 3904
rect 1610 3524 1622 3526
rect 1610 3516 1612 3524
rect 1620 3516 1622 3524
rect 1610 3304 1622 3516
rect 1610 3296 1612 3304
rect 1620 3296 1622 3304
rect 1610 3294 1622 3296
rect 1674 2964 1686 3896
rect 1930 3584 1942 3586
rect 1930 3576 1932 3584
rect 1940 3576 1942 3584
rect 1674 2956 1676 2964
rect 1684 2956 1686 2964
rect 1674 2954 1686 2956
rect 1706 3484 1718 3486
rect 1706 3476 1708 3484
rect 1716 3476 1718 3484
rect 1706 3444 1718 3476
rect 1706 3436 1708 3444
rect 1716 3436 1718 3444
rect 1578 2776 1580 2784
rect 1588 2776 1590 2784
rect 1578 2774 1590 2776
rect 1706 2744 1718 3436
rect 1898 3404 1910 3406
rect 1898 3396 1900 3404
rect 1908 3396 1910 3404
rect 1866 3324 1878 3326
rect 1866 3316 1868 3324
rect 1876 3316 1878 3324
rect 1834 3304 1846 3306
rect 1834 3296 1836 3304
rect 1844 3296 1846 3304
rect 1834 3124 1846 3296
rect 1834 3116 1836 3124
rect 1844 3116 1846 3124
rect 1834 3114 1846 3116
rect 1866 2924 1878 3316
rect 1866 2916 1868 2924
rect 1876 2916 1878 2924
rect 1866 2914 1878 2916
rect 1834 2904 1846 2906
rect 1834 2896 1836 2904
rect 1844 2896 1846 2904
rect 1706 2736 1708 2744
rect 1716 2736 1718 2744
rect 1706 2734 1718 2736
rect 1770 2824 1782 2826
rect 1770 2816 1772 2824
rect 1780 2816 1782 2824
rect 1578 2704 1590 2706
rect 1578 2696 1580 2704
rect 1588 2696 1590 2704
rect 1578 2444 1590 2696
rect 1674 2704 1686 2706
rect 1674 2696 1676 2704
rect 1684 2696 1686 2704
rect 1674 2664 1686 2696
rect 1674 2656 1676 2664
rect 1684 2656 1686 2664
rect 1674 2654 1686 2656
rect 1578 2436 1580 2444
rect 1588 2436 1590 2444
rect 1578 2434 1590 2436
rect 1738 2424 1750 2426
rect 1738 2416 1740 2424
rect 1748 2416 1750 2424
rect 1706 1924 1718 1926
rect 1706 1916 1708 1924
rect 1716 1916 1718 1924
rect 1642 1784 1654 1786
rect 1642 1776 1644 1784
rect 1652 1776 1654 1784
rect 1642 1724 1654 1776
rect 1642 1716 1644 1724
rect 1652 1716 1654 1724
rect 1642 1714 1654 1716
rect 1674 1724 1686 1726
rect 1674 1716 1676 1724
rect 1684 1716 1686 1724
rect 1514 1616 1516 1624
rect 1524 1616 1526 1624
rect 1514 1614 1526 1616
rect 1610 1624 1622 1626
rect 1610 1616 1612 1624
rect 1620 1616 1622 1624
rect 1408 1606 1412 1614
rect 1420 1606 1424 1614
rect 1432 1606 1436 1614
rect 1444 1606 1448 1614
rect 1456 1606 1460 1614
rect 1468 1606 1472 1614
rect 1258 1456 1260 1464
rect 1268 1456 1270 1464
rect 1258 1454 1270 1456
rect 1354 1544 1366 1546
rect 1354 1536 1356 1544
rect 1364 1536 1366 1544
rect 1226 1396 1228 1404
rect 1236 1396 1238 1404
rect 1226 1394 1238 1396
rect 1258 1404 1270 1406
rect 1258 1396 1260 1404
rect 1268 1396 1270 1404
rect 1098 996 1100 1004
rect 1108 996 1110 1004
rect 1098 994 1110 996
rect 1258 844 1270 1396
rect 1322 1244 1334 1246
rect 1322 1236 1324 1244
rect 1332 1236 1334 1244
rect 1290 944 1302 946
rect 1290 936 1292 944
rect 1300 936 1302 944
rect 1290 884 1302 936
rect 1290 876 1292 884
rect 1300 876 1302 884
rect 1290 874 1302 876
rect 1258 836 1260 844
rect 1268 836 1270 844
rect 1258 834 1270 836
rect 1002 676 1004 684
rect 1012 676 1014 684
rect 1002 674 1014 676
rect 1034 764 1046 766
rect 1034 756 1036 764
rect 1044 756 1046 764
rect 778 296 780 304
rect 788 296 790 304
rect 778 294 790 296
rect 810 644 822 646
rect 810 636 812 644
rect 820 636 822 644
rect 362 156 364 164
rect 372 156 374 164
rect 362 154 374 156
rect 810 164 822 636
rect 842 284 886 286
rect 842 276 844 284
rect 852 276 886 284
rect 842 274 886 276
rect 874 264 886 274
rect 874 256 876 264
rect 884 256 886 264
rect 874 254 886 256
rect 1034 184 1046 756
rect 1162 724 1174 726
rect 1162 716 1164 724
rect 1172 716 1174 724
rect 1162 564 1174 716
rect 1162 556 1164 564
rect 1172 556 1174 564
rect 1162 304 1174 556
rect 1322 504 1334 1236
rect 1354 1084 1366 1536
rect 1354 1076 1356 1084
rect 1364 1076 1366 1084
rect 1354 1074 1366 1076
rect 1408 1214 1472 1606
rect 1546 1504 1558 1506
rect 1546 1496 1548 1504
rect 1556 1496 1558 1504
rect 1546 1304 1558 1496
rect 1546 1296 1548 1304
rect 1556 1296 1558 1304
rect 1546 1294 1558 1296
rect 1578 1444 1590 1446
rect 1578 1436 1580 1444
rect 1588 1436 1590 1444
rect 1408 1206 1412 1214
rect 1420 1206 1424 1214
rect 1432 1206 1436 1214
rect 1444 1206 1448 1214
rect 1456 1206 1460 1214
rect 1468 1206 1472 1214
rect 1322 496 1324 504
rect 1332 496 1334 504
rect 1322 494 1334 496
rect 1408 814 1472 1206
rect 1578 1204 1590 1436
rect 1578 1196 1580 1204
rect 1588 1196 1590 1204
rect 1578 1194 1590 1196
rect 1610 884 1622 1616
rect 1674 1444 1686 1716
rect 1706 1644 1718 1916
rect 1706 1636 1708 1644
rect 1716 1636 1718 1644
rect 1706 1634 1718 1636
rect 1674 1436 1676 1444
rect 1684 1436 1686 1444
rect 1674 1434 1686 1436
rect 1706 1444 1718 1446
rect 1706 1436 1708 1444
rect 1716 1436 1718 1444
rect 1706 1224 1718 1436
rect 1706 1216 1708 1224
rect 1716 1216 1718 1224
rect 1706 1214 1718 1216
rect 1674 1164 1686 1166
rect 1674 1156 1676 1164
rect 1684 1156 1686 1164
rect 1674 1064 1686 1156
rect 1674 1056 1676 1064
rect 1684 1056 1686 1064
rect 1674 1054 1686 1056
rect 1610 876 1612 884
rect 1620 876 1622 884
rect 1610 874 1622 876
rect 1408 806 1412 814
rect 1420 806 1424 814
rect 1432 806 1436 814
rect 1444 806 1448 814
rect 1456 806 1460 814
rect 1468 806 1472 814
rect 1162 296 1164 304
rect 1172 296 1174 304
rect 1162 294 1174 296
rect 1408 414 1472 806
rect 1738 504 1750 2416
rect 1770 2424 1782 2816
rect 1770 2416 1772 2424
rect 1780 2416 1782 2424
rect 1770 2414 1782 2416
rect 1802 2824 1814 2826
rect 1802 2816 1804 2824
rect 1812 2816 1814 2824
rect 1802 2344 1814 2816
rect 1802 2336 1804 2344
rect 1812 2336 1814 2344
rect 1802 2334 1814 2336
rect 1834 2284 1846 2896
rect 1898 2764 1910 3396
rect 1930 3164 1942 3576
rect 2058 3504 2070 3506
rect 2058 3496 2060 3504
rect 2068 3496 2070 3504
rect 1930 3156 1932 3164
rect 1940 3156 1942 3164
rect 1930 3154 1942 3156
rect 1962 3484 1974 3486
rect 1962 3476 1964 3484
rect 1972 3476 1974 3484
rect 1898 2756 1900 2764
rect 1908 2756 1910 2764
rect 1898 2754 1910 2756
rect 1962 2664 1974 3476
rect 2058 2904 2070 3496
rect 2058 2896 2060 2904
rect 2068 2896 2070 2904
rect 2058 2894 2070 2896
rect 1962 2656 1964 2664
rect 1972 2656 1974 2664
rect 1962 2654 1974 2656
rect 1898 2644 1910 2646
rect 1898 2636 1900 2644
rect 1908 2636 1910 2644
rect 1898 2424 1910 2636
rect 1994 2524 2006 2526
rect 1994 2516 1996 2524
rect 2004 2516 2006 2524
rect 1994 2464 2006 2516
rect 2122 2484 2134 4296
rect 2250 4244 2262 4936
rect 2378 4944 2390 4946
rect 2378 4936 2380 4944
rect 2388 4936 2390 4944
rect 2250 4236 2252 4244
rect 2260 4236 2262 4244
rect 2250 4234 2262 4236
rect 2282 4704 2294 4706
rect 2282 4696 2284 4704
rect 2292 4696 2294 4704
rect 2218 4204 2230 4206
rect 2218 4196 2220 4204
rect 2228 4196 2230 4204
rect 2154 3164 2166 3166
rect 2154 3156 2156 3164
rect 2164 3156 2166 3164
rect 2154 2844 2166 3156
rect 2154 2836 2156 2844
rect 2164 2836 2166 2844
rect 2154 2834 2166 2836
rect 2218 2644 2230 4196
rect 2282 4104 2294 4696
rect 2378 4564 2390 4936
rect 2410 4844 2422 4976
rect 2410 4836 2412 4844
rect 2420 4836 2422 4844
rect 2410 4834 2422 4836
rect 2570 4764 2582 5016
rect 2570 4756 2572 4764
rect 2580 4756 2582 4764
rect 2570 4754 2582 4756
rect 2602 4784 2614 4786
rect 2602 4776 2604 4784
rect 2612 4776 2614 4784
rect 2378 4556 2380 4564
rect 2388 4556 2390 4564
rect 2378 4554 2390 4556
rect 2570 4544 2582 4546
rect 2570 4536 2572 4544
rect 2580 4536 2582 4544
rect 2570 4144 2582 4536
rect 2602 4544 2614 4776
rect 2602 4536 2604 4544
rect 2612 4536 2614 4544
rect 2602 4534 2614 4536
rect 2570 4136 2572 4144
rect 2580 4136 2582 4144
rect 2570 4134 2582 4136
rect 2282 4096 2284 4104
rect 2292 4096 2294 4104
rect 2282 4094 2294 4096
rect 2410 4084 2422 4086
rect 2410 4076 2412 4084
rect 2420 4076 2422 4084
rect 2314 3744 2326 3746
rect 2314 3736 2316 3744
rect 2324 3736 2326 3744
rect 2314 3484 2326 3736
rect 2314 3476 2316 3484
rect 2324 3476 2326 3484
rect 2314 3474 2326 3476
rect 2346 3204 2358 3206
rect 2346 3196 2348 3204
rect 2356 3196 2358 3204
rect 2218 2636 2220 2644
rect 2228 2636 2230 2644
rect 2218 2634 2230 2636
rect 2250 2744 2262 2746
rect 2250 2736 2252 2744
rect 2260 2736 2262 2744
rect 2186 2504 2198 2506
rect 2186 2496 2188 2504
rect 2196 2496 2198 2504
rect 2122 2476 2124 2484
rect 2132 2476 2134 2484
rect 2122 2474 2134 2476
rect 2154 2484 2166 2486
rect 2154 2476 2156 2484
rect 2164 2476 2166 2484
rect 1994 2456 1996 2464
rect 2004 2456 2006 2464
rect 1994 2454 2006 2456
rect 1898 2416 1900 2424
rect 1908 2416 1910 2424
rect 1898 2414 1910 2416
rect 1834 2276 1836 2284
rect 1844 2276 1846 2284
rect 1834 1744 1846 2276
rect 1962 2344 1974 2346
rect 1962 2336 1964 2344
rect 1972 2336 1974 2344
rect 1962 2144 1974 2336
rect 1962 2136 1964 2144
rect 1972 2136 1974 2144
rect 1866 2104 1878 2106
rect 1866 2096 1868 2104
rect 1876 2096 1878 2104
rect 1866 2024 1878 2096
rect 1866 2016 1868 2024
rect 1876 2016 1878 2024
rect 1866 2014 1878 2016
rect 1834 1736 1836 1744
rect 1844 1736 1846 1744
rect 1834 1734 1846 1736
rect 1962 1844 1974 2136
rect 1962 1836 1964 1844
rect 1972 1836 1974 1844
rect 1962 1724 1974 1836
rect 1962 1716 1964 1724
rect 1972 1716 1974 1724
rect 1962 1714 1974 1716
rect 1994 2324 2006 2326
rect 1994 2316 1996 2324
rect 2004 2316 2006 2324
rect 1994 1724 2006 2316
rect 2090 2304 2102 2306
rect 2090 2296 2092 2304
rect 2100 2296 2102 2304
rect 2090 2164 2102 2296
rect 2090 2156 2092 2164
rect 2100 2156 2102 2164
rect 2090 2154 2102 2156
rect 1994 1716 1996 1724
rect 2004 1716 2006 1724
rect 1994 1714 2006 1716
rect 2154 1684 2166 2476
rect 2186 2184 2198 2496
rect 2186 2176 2188 2184
rect 2196 2176 2198 2184
rect 2186 2174 2198 2176
rect 2250 2324 2262 2736
rect 2250 2316 2252 2324
rect 2260 2316 2262 2324
rect 2250 2104 2262 2316
rect 2250 2096 2252 2104
rect 2260 2096 2262 2104
rect 2250 2094 2262 2096
rect 2282 2644 2294 2646
rect 2282 2636 2284 2644
rect 2292 2636 2294 2644
rect 2186 1944 2198 1946
rect 2186 1936 2188 1944
rect 2196 1936 2198 1944
rect 2186 1864 2198 1936
rect 2186 1856 2188 1864
rect 2196 1856 2198 1864
rect 2186 1854 2198 1856
rect 2250 1884 2262 1886
rect 2250 1876 2252 1884
rect 2260 1876 2262 1884
rect 2154 1676 2156 1684
rect 2164 1676 2166 1684
rect 2154 1674 2166 1676
rect 2218 1824 2230 1826
rect 2218 1816 2220 1824
rect 2228 1816 2230 1824
rect 2218 1684 2230 1816
rect 2250 1704 2262 1876
rect 2282 1724 2294 2636
rect 2314 2064 2326 2066
rect 2314 2056 2316 2064
rect 2324 2056 2326 2064
rect 2314 2004 2326 2056
rect 2314 1996 2316 2004
rect 2324 1996 2326 2004
rect 2314 1994 2326 1996
rect 2346 1884 2358 3196
rect 2410 3104 2422 4076
rect 2474 3904 2486 3906
rect 2474 3896 2476 3904
rect 2484 3896 2486 3904
rect 2474 3724 2486 3896
rect 2570 3904 2582 3906
rect 2570 3896 2572 3904
rect 2580 3896 2582 3904
rect 2474 3716 2476 3724
rect 2484 3716 2486 3724
rect 2474 3714 2486 3716
rect 2506 3804 2518 3806
rect 2506 3796 2508 3804
rect 2516 3796 2518 3804
rect 2410 3096 2412 3104
rect 2420 3096 2422 3104
rect 2410 3094 2422 3096
rect 2474 3524 2486 3526
rect 2474 3516 2476 3524
rect 2484 3516 2486 3524
rect 2378 3004 2390 3006
rect 2378 2996 2380 3004
rect 2388 2996 2390 3004
rect 2378 2924 2390 2996
rect 2378 2916 2380 2924
rect 2388 2916 2390 2924
rect 2378 2914 2390 2916
rect 2474 2884 2486 3516
rect 2506 3484 2518 3796
rect 2570 3544 2582 3896
rect 2634 3884 2646 3886
rect 2634 3876 2636 3884
rect 2644 3876 2646 3884
rect 2634 3724 2646 3876
rect 2634 3716 2636 3724
rect 2644 3716 2646 3724
rect 2634 3714 2646 3716
rect 2666 3644 2678 5176
rect 2912 5014 2976 5406
rect 2912 5006 2916 5014
rect 2924 5006 2928 5014
rect 2936 5006 2940 5014
rect 2948 5006 2952 5014
rect 2960 5006 2964 5014
rect 2972 5006 2976 5014
rect 2912 4614 2976 5006
rect 3210 5304 3222 5306
rect 3210 5296 3212 5304
rect 3220 5296 3222 5304
rect 2912 4606 2916 4614
rect 2924 4606 2928 4614
rect 2936 4606 2940 4614
rect 2948 4606 2952 4614
rect 2960 4606 2964 4614
rect 2972 4606 2976 4614
rect 2762 4564 2774 4566
rect 2762 4556 2764 4564
rect 2772 4556 2774 4564
rect 2762 4084 2774 4556
rect 2762 4076 2764 4084
rect 2772 4076 2774 4084
rect 2762 4074 2774 4076
rect 2794 4444 2806 4446
rect 2794 4436 2796 4444
rect 2804 4436 2806 4444
rect 2666 3636 2668 3644
rect 2676 3636 2678 3644
rect 2666 3634 2678 3636
rect 2730 4044 2742 4046
rect 2730 4036 2732 4044
rect 2740 4036 2742 4044
rect 2570 3536 2572 3544
rect 2580 3536 2582 3544
rect 2570 3534 2582 3536
rect 2506 3476 2508 3484
rect 2516 3476 2518 3484
rect 2506 3474 2518 3476
rect 2698 3504 2710 3506
rect 2698 3496 2700 3504
rect 2708 3496 2710 3504
rect 2698 3364 2710 3496
rect 2730 3484 2742 4036
rect 2730 3476 2732 3484
rect 2740 3476 2742 3484
rect 2730 3474 2742 3476
rect 2698 3356 2700 3364
rect 2708 3356 2710 3364
rect 2698 3354 2710 3356
rect 2474 2876 2476 2884
rect 2484 2876 2486 2884
rect 2474 2874 2486 2876
rect 2570 3124 2582 3126
rect 2570 3116 2572 3124
rect 2580 3116 2582 3124
rect 2442 2864 2454 2866
rect 2442 2856 2444 2864
rect 2452 2856 2454 2864
rect 2378 2824 2390 2826
rect 2378 2816 2380 2824
rect 2388 2816 2390 2824
rect 2378 2064 2390 2816
rect 2410 2684 2422 2686
rect 2410 2676 2412 2684
rect 2420 2676 2422 2684
rect 2410 2444 2422 2676
rect 2410 2436 2412 2444
rect 2420 2436 2422 2444
rect 2410 2434 2422 2436
rect 2442 2304 2454 2856
rect 2442 2296 2444 2304
rect 2452 2296 2454 2304
rect 2442 2294 2454 2296
rect 2474 2684 2486 2686
rect 2474 2676 2476 2684
rect 2484 2676 2486 2684
rect 2378 2056 2380 2064
rect 2388 2056 2390 2064
rect 2378 2054 2390 2056
rect 2346 1876 2348 1884
rect 2356 1876 2358 1884
rect 2346 1874 2358 1876
rect 2378 1904 2390 1906
rect 2378 1896 2380 1904
rect 2388 1896 2390 1904
rect 2314 1844 2326 1846
rect 2314 1836 2316 1844
rect 2324 1836 2326 1844
rect 2314 1784 2326 1836
rect 2314 1776 2316 1784
rect 2324 1776 2326 1784
rect 2314 1774 2326 1776
rect 2346 1844 2358 1846
rect 2346 1836 2348 1844
rect 2356 1836 2358 1844
rect 2282 1716 2284 1724
rect 2292 1716 2294 1724
rect 2282 1714 2294 1716
rect 2250 1696 2252 1704
rect 2260 1696 2262 1704
rect 2250 1694 2262 1696
rect 2218 1676 2220 1684
rect 2228 1676 2230 1684
rect 2218 1674 2230 1676
rect 2186 1524 2198 1526
rect 2186 1516 2188 1524
rect 2196 1516 2198 1524
rect 1898 1224 1910 1226
rect 1898 1216 1900 1224
rect 1908 1216 1910 1224
rect 1898 884 1910 1216
rect 2122 1064 2134 1066
rect 2122 1056 2124 1064
rect 2132 1056 2134 1064
rect 2090 984 2102 986
rect 2090 976 2092 984
rect 2100 976 2102 984
rect 1898 876 1900 884
rect 1908 876 1910 884
rect 1898 874 1910 876
rect 2058 924 2070 926
rect 2058 916 2060 924
rect 2068 916 2070 924
rect 2058 884 2070 916
rect 2090 924 2102 976
rect 2090 916 2092 924
rect 2100 916 2102 924
rect 2090 914 2102 916
rect 2058 876 2060 884
rect 2068 876 2070 884
rect 2058 874 2070 876
rect 2122 884 2134 1056
rect 2122 876 2124 884
rect 2132 876 2134 884
rect 2122 874 2134 876
rect 1866 784 1878 786
rect 1866 776 1868 784
rect 1876 776 1878 784
rect 1866 524 1878 776
rect 2154 684 2166 686
rect 2154 676 2156 684
rect 2164 676 2166 684
rect 2154 544 2166 676
rect 2154 536 2156 544
rect 2164 536 2166 544
rect 2154 534 2166 536
rect 1866 516 1868 524
rect 1876 516 1878 524
rect 1866 514 1878 516
rect 1738 496 1740 504
rect 1748 496 1750 504
rect 1738 494 1750 496
rect 2186 504 2198 1516
rect 2346 1264 2358 1836
rect 2378 1724 2390 1896
rect 2378 1716 2380 1724
rect 2388 1716 2390 1724
rect 2378 1714 2390 1716
rect 2410 1484 2422 1486
rect 2410 1476 2412 1484
rect 2420 1476 2422 1484
rect 2410 1324 2422 1476
rect 2410 1316 2412 1324
rect 2420 1316 2422 1324
rect 2410 1314 2422 1316
rect 2346 1256 2348 1264
rect 2356 1256 2358 1264
rect 2346 1254 2358 1256
rect 2474 1204 2486 2676
rect 2506 2284 2518 2286
rect 2506 2276 2508 2284
rect 2516 2276 2518 2284
rect 2506 2064 2518 2276
rect 2570 2264 2582 3116
rect 2698 3004 2710 3006
rect 2698 2996 2700 3004
rect 2708 2996 2710 3004
rect 2634 2824 2646 2826
rect 2634 2816 2636 2824
rect 2644 2816 2646 2824
rect 2570 2256 2572 2264
rect 2580 2256 2582 2264
rect 2570 2254 2582 2256
rect 2602 2424 2614 2426
rect 2602 2416 2604 2424
rect 2612 2416 2614 2424
rect 2602 2264 2614 2416
rect 2602 2256 2604 2264
rect 2612 2256 2614 2264
rect 2602 2254 2614 2256
rect 2570 2144 2582 2146
rect 2570 2136 2572 2144
rect 2580 2136 2582 2144
rect 2506 2056 2508 2064
rect 2516 2056 2518 2064
rect 2506 2054 2518 2056
rect 2538 2104 2550 2106
rect 2538 2096 2540 2104
rect 2548 2096 2550 2104
rect 2538 1444 2550 2096
rect 2570 1864 2582 2136
rect 2634 2104 2646 2816
rect 2698 2764 2710 2996
rect 2698 2756 2700 2764
rect 2708 2756 2710 2764
rect 2698 2754 2710 2756
rect 2698 2724 2710 2726
rect 2698 2716 2700 2724
rect 2708 2716 2710 2724
rect 2698 2524 2710 2716
rect 2698 2516 2700 2524
rect 2708 2516 2710 2524
rect 2698 2514 2710 2516
rect 2762 2684 2774 2686
rect 2762 2676 2764 2684
rect 2772 2676 2774 2684
rect 2762 2284 2774 2676
rect 2794 2524 2806 4436
rect 2912 4214 2976 4606
rect 3082 4964 3094 4966
rect 3082 4956 3084 4964
rect 3092 4956 3094 4964
rect 3082 4544 3094 4956
rect 3210 4844 3222 5296
rect 3434 5284 3446 5416
rect 3434 5276 3436 5284
rect 3444 5276 3446 5284
rect 3434 5274 3446 5276
rect 3466 5424 3478 5426
rect 3466 5416 3468 5424
rect 3476 5416 3478 5424
rect 3434 5164 3446 5166
rect 3434 5156 3436 5164
rect 3444 5156 3446 5164
rect 3434 5064 3446 5156
rect 3434 5056 3436 5064
rect 3444 5056 3446 5064
rect 3434 5054 3446 5056
rect 3210 4836 3212 4844
rect 3220 4836 3222 4844
rect 3210 4834 3222 4836
rect 3402 4944 3414 4946
rect 3402 4936 3404 4944
rect 3412 4936 3414 4944
rect 3338 4824 3350 4826
rect 3338 4816 3340 4824
rect 3348 4816 3350 4824
rect 3082 4536 3084 4544
rect 3092 4536 3094 4544
rect 3082 4534 3094 4536
rect 3146 4704 3158 4706
rect 3146 4696 3148 4704
rect 3156 4696 3158 4704
rect 2912 4206 2916 4214
rect 2924 4206 2928 4214
rect 2936 4206 2940 4214
rect 2948 4206 2952 4214
rect 2960 4206 2964 4214
rect 2972 4206 2976 4214
rect 2912 3814 2976 4206
rect 3082 4224 3094 4226
rect 3082 4216 3084 4224
rect 3092 4216 3094 4224
rect 3082 4084 3094 4216
rect 3082 4076 3084 4084
rect 3092 4076 3094 4084
rect 3082 4074 3094 4076
rect 2912 3806 2916 3814
rect 2924 3806 2928 3814
rect 2936 3806 2940 3814
rect 2948 3806 2952 3814
rect 2960 3806 2964 3814
rect 2972 3806 2976 3814
rect 2912 3414 2976 3806
rect 2912 3406 2916 3414
rect 2924 3406 2928 3414
rect 2936 3406 2940 3414
rect 2948 3406 2952 3414
rect 2960 3406 2964 3414
rect 2972 3406 2976 3414
rect 2912 3014 2976 3406
rect 3114 4064 3126 4066
rect 3114 4056 3116 4064
rect 3124 4056 3126 4064
rect 3114 3364 3126 4056
rect 3146 4024 3158 4696
rect 3242 4444 3254 4446
rect 3242 4436 3244 4444
rect 3252 4436 3254 4444
rect 3242 4104 3254 4436
rect 3242 4096 3244 4104
rect 3252 4096 3254 4104
rect 3242 4094 3254 4096
rect 3274 4424 3286 4426
rect 3274 4416 3276 4424
rect 3284 4416 3286 4424
rect 3146 4016 3148 4024
rect 3156 4016 3158 4024
rect 3146 4014 3158 4016
rect 3114 3356 3116 3364
rect 3124 3356 3126 3364
rect 3114 3354 3126 3356
rect 3146 3984 3158 3986
rect 3146 3976 3148 3984
rect 3156 3976 3158 3984
rect 2912 3006 2916 3014
rect 2924 3006 2928 3014
rect 2936 3006 2940 3014
rect 2948 3006 2952 3014
rect 2960 3006 2964 3014
rect 2972 3006 2976 3014
rect 2912 2614 2976 3006
rect 2912 2606 2916 2614
rect 2924 2606 2928 2614
rect 2936 2606 2940 2614
rect 2948 2606 2952 2614
rect 2960 2606 2964 2614
rect 2972 2606 2976 2614
rect 2794 2516 2796 2524
rect 2804 2516 2806 2524
rect 2794 2514 2806 2516
rect 2858 2544 2870 2546
rect 2858 2536 2860 2544
rect 2868 2536 2870 2544
rect 2762 2276 2764 2284
rect 2772 2276 2774 2284
rect 2762 2274 2774 2276
rect 2634 2096 2636 2104
rect 2644 2096 2646 2104
rect 2634 2094 2646 2096
rect 2666 2264 2678 2266
rect 2666 2256 2668 2264
rect 2676 2256 2678 2264
rect 2634 1944 2646 1946
rect 2634 1936 2636 1944
rect 2644 1936 2646 1944
rect 2570 1856 2572 1864
rect 2580 1856 2582 1864
rect 2570 1854 2582 1856
rect 2602 1864 2614 1866
rect 2602 1856 2604 1864
rect 2612 1856 2614 1864
rect 2570 1744 2582 1746
rect 2570 1736 2572 1744
rect 2580 1736 2582 1744
rect 2570 1644 2582 1736
rect 2570 1636 2572 1644
rect 2580 1636 2582 1644
rect 2570 1634 2582 1636
rect 2538 1436 2540 1444
rect 2548 1436 2550 1444
rect 2538 1434 2550 1436
rect 2506 1344 2518 1346
rect 2506 1336 2508 1344
rect 2516 1336 2518 1344
rect 2506 1304 2518 1336
rect 2602 1344 2614 1856
rect 2634 1804 2646 1936
rect 2634 1796 2636 1804
rect 2644 1796 2646 1804
rect 2634 1794 2646 1796
rect 2666 1664 2678 2256
rect 2666 1656 2668 1664
rect 2676 1656 2678 1664
rect 2666 1654 2678 1656
rect 2698 2264 2710 2266
rect 2698 2256 2700 2264
rect 2708 2256 2710 2264
rect 2698 1644 2710 2256
rect 2858 2244 2870 2536
rect 2858 2236 2860 2244
rect 2868 2236 2870 2244
rect 2858 2234 2870 2236
rect 2730 2224 2742 2226
rect 2730 2216 2732 2224
rect 2740 2216 2742 2224
rect 2730 2104 2742 2216
rect 2912 2214 2976 2606
rect 3114 3304 3126 3306
rect 3114 3296 3116 3304
rect 3124 3296 3126 3304
rect 3082 2344 3094 2346
rect 3082 2336 3084 2344
rect 3092 2336 3094 2344
rect 2912 2206 2916 2214
rect 2924 2206 2928 2214
rect 2936 2206 2940 2214
rect 2948 2206 2952 2214
rect 2960 2206 2964 2214
rect 2972 2206 2976 2214
rect 2730 2096 2732 2104
rect 2740 2096 2742 2104
rect 2730 2094 2742 2096
rect 2794 2204 2806 2206
rect 2794 2196 2796 2204
rect 2804 2196 2806 2204
rect 2794 2104 2806 2196
rect 2794 2096 2796 2104
rect 2804 2096 2806 2104
rect 2794 2094 2806 2096
rect 2826 2124 2838 2126
rect 2826 2116 2828 2124
rect 2836 2116 2838 2124
rect 2698 1636 2700 1644
rect 2708 1636 2710 1644
rect 2698 1634 2710 1636
rect 2730 2064 2742 2066
rect 2730 2056 2732 2064
rect 2740 2056 2742 2064
rect 2730 1584 2742 2056
rect 2730 1576 2732 1584
rect 2740 1576 2742 1584
rect 2730 1574 2742 1576
rect 2762 2064 2774 2066
rect 2762 2056 2764 2064
rect 2772 2056 2774 2064
rect 2762 1464 2774 2056
rect 2826 1864 2838 2116
rect 2826 1856 2828 1864
rect 2836 1856 2838 1864
rect 2826 1854 2838 1856
rect 2762 1456 2764 1464
rect 2772 1456 2774 1464
rect 2762 1454 2774 1456
rect 2912 1814 2976 2206
rect 3018 2284 3030 2286
rect 3018 2276 3020 2284
rect 3028 2276 3030 2284
rect 3018 2124 3030 2276
rect 3018 2116 3020 2124
rect 3028 2116 3030 2124
rect 3018 2114 3030 2116
rect 2912 1806 2916 1814
rect 2924 1806 2928 1814
rect 2936 1806 2940 1814
rect 2948 1806 2952 1814
rect 2960 1806 2964 1814
rect 2972 1806 2976 1814
rect 2602 1336 2604 1344
rect 2612 1336 2614 1344
rect 2602 1334 2614 1336
rect 2912 1414 2976 1806
rect 2912 1406 2916 1414
rect 2924 1406 2928 1414
rect 2936 1406 2940 1414
rect 2948 1406 2952 1414
rect 2960 1406 2964 1414
rect 2972 1406 2976 1414
rect 2506 1296 2508 1304
rect 2516 1296 2518 1304
rect 2506 1294 2518 1296
rect 2474 1196 2476 1204
rect 2484 1196 2486 1204
rect 2474 1194 2486 1196
rect 2858 1124 2870 1126
rect 2858 1116 2860 1124
rect 2868 1116 2870 1124
rect 2314 1104 2326 1106
rect 2314 1096 2316 1104
rect 2324 1096 2326 1104
rect 2218 984 2230 986
rect 2218 976 2220 984
rect 2228 976 2230 984
rect 2218 924 2230 976
rect 2218 916 2220 924
rect 2228 916 2230 924
rect 2218 914 2230 916
rect 2314 744 2326 1096
rect 2538 1064 2550 1066
rect 2538 1056 2540 1064
rect 2548 1056 2550 1064
rect 2314 736 2316 744
rect 2324 736 2326 744
rect 2314 734 2326 736
rect 2442 764 2454 766
rect 2442 756 2444 764
rect 2452 756 2454 764
rect 2282 704 2294 706
rect 2282 696 2284 704
rect 2292 696 2294 704
rect 2282 664 2294 696
rect 2282 656 2284 664
rect 2292 656 2294 664
rect 2282 654 2294 656
rect 2186 496 2188 504
rect 2196 496 2198 504
rect 2186 494 2198 496
rect 2442 484 2454 756
rect 2538 664 2550 1056
rect 2538 656 2540 664
rect 2548 656 2550 664
rect 2538 654 2550 656
rect 2570 864 2582 866
rect 2570 856 2572 864
rect 2580 856 2582 864
rect 2474 624 2486 626
rect 2474 616 2476 624
rect 2484 616 2486 624
rect 2474 584 2486 616
rect 2474 576 2476 584
rect 2484 576 2486 584
rect 2474 574 2486 576
rect 2442 476 2444 484
rect 2452 476 2454 484
rect 2442 474 2454 476
rect 2570 484 2582 856
rect 2858 724 2870 1116
rect 2858 716 2860 724
rect 2868 716 2870 724
rect 2858 714 2870 716
rect 2912 1014 2976 1406
rect 3018 1624 3030 1626
rect 3018 1616 3020 1624
rect 3028 1616 3030 1624
rect 3018 1024 3030 1616
rect 3050 1624 3062 1626
rect 3050 1616 3052 1624
rect 3060 1616 3062 1624
rect 3050 1344 3062 1616
rect 3082 1404 3094 2336
rect 3082 1396 3084 1404
rect 3092 1396 3094 1404
rect 3082 1394 3094 1396
rect 3114 2324 3126 3296
rect 3146 2584 3158 3976
rect 3274 3964 3286 4416
rect 3338 4244 3350 4816
rect 3338 4236 3340 4244
rect 3348 4236 3350 4244
rect 3338 4234 3350 4236
rect 3370 4204 3382 4206
rect 3370 4196 3372 4204
rect 3380 4196 3382 4204
rect 3274 3956 3276 3964
rect 3284 3956 3286 3964
rect 3274 3954 3286 3956
rect 3306 3984 3318 3986
rect 3306 3976 3308 3984
rect 3316 3976 3318 3984
rect 3306 2884 3318 3976
rect 3338 3724 3350 3726
rect 3338 3716 3340 3724
rect 3348 3716 3350 3724
rect 3338 3264 3350 3716
rect 3370 3604 3382 4196
rect 3402 4204 3414 4936
rect 3466 4904 3478 5416
rect 3562 5404 3574 5406
rect 3562 5396 3564 5404
rect 3572 5396 3574 5404
rect 3466 4896 3468 4904
rect 3476 4896 3478 4904
rect 3466 4894 3478 4896
rect 3530 5104 3542 5106
rect 3530 5096 3532 5104
rect 3540 5096 3542 5104
rect 3466 4844 3478 4846
rect 3466 4836 3468 4844
rect 3476 4836 3478 4844
rect 3402 4196 3404 4204
rect 3412 4196 3414 4204
rect 3402 4194 3414 4196
rect 3434 4604 3446 4606
rect 3434 4596 3436 4604
rect 3444 4596 3446 4604
rect 3370 3596 3372 3604
rect 3380 3596 3382 3604
rect 3370 3594 3382 3596
rect 3402 4144 3414 4146
rect 3402 4136 3404 4144
rect 3412 4136 3414 4144
rect 3402 3484 3414 4136
rect 3434 3584 3446 4596
rect 3466 4504 3478 4836
rect 3466 4496 3468 4504
rect 3476 4496 3478 4504
rect 3466 4494 3478 4496
rect 3498 4784 3510 4786
rect 3498 4776 3500 4784
rect 3508 4776 3510 4784
rect 3498 4444 3510 4776
rect 3498 4436 3500 4444
rect 3508 4436 3510 4444
rect 3498 4434 3510 4436
rect 3530 4504 3542 5096
rect 3562 4564 3574 5396
rect 4010 5304 4022 5306
rect 4010 5296 4012 5304
rect 4020 5296 4022 5304
rect 3786 4964 3798 4966
rect 3786 4956 3788 4964
rect 3796 4956 3798 4964
rect 3626 4804 3638 4806
rect 3626 4796 3628 4804
rect 3636 4796 3638 4804
rect 3562 4556 3564 4564
rect 3572 4556 3574 4564
rect 3562 4554 3574 4556
rect 3594 4704 3606 4706
rect 3594 4696 3596 4704
rect 3604 4696 3606 4704
rect 3530 4496 3532 4504
rect 3540 4496 3542 4504
rect 3498 4404 3510 4406
rect 3498 4396 3500 4404
rect 3508 4396 3510 4404
rect 3498 4244 3510 4396
rect 3498 4236 3500 4244
rect 3508 4236 3510 4244
rect 3498 4234 3510 4236
rect 3466 4164 3478 4166
rect 3466 4156 3468 4164
rect 3476 4156 3478 4164
rect 3466 4004 3478 4156
rect 3466 3996 3468 4004
rect 3476 3996 3478 4004
rect 3466 3994 3478 3996
rect 3434 3576 3436 3584
rect 3444 3576 3446 3584
rect 3434 3574 3446 3576
rect 3402 3476 3404 3484
rect 3412 3476 3414 3484
rect 3402 3474 3414 3476
rect 3338 3256 3340 3264
rect 3348 3256 3350 3264
rect 3338 3254 3350 3256
rect 3466 2904 3478 2906
rect 3466 2896 3468 2904
rect 3476 2896 3478 2904
rect 3306 2876 3308 2884
rect 3316 2876 3318 2884
rect 3306 2874 3318 2876
rect 3370 2884 3382 2886
rect 3370 2876 3372 2884
rect 3380 2876 3382 2884
rect 3146 2576 3148 2584
rect 3156 2576 3158 2584
rect 3146 2574 3158 2576
rect 3114 2316 3116 2324
rect 3124 2316 3126 2324
rect 3114 2104 3126 2316
rect 3114 2096 3116 2104
rect 3124 2096 3126 2104
rect 3050 1336 3052 1344
rect 3060 1336 3062 1344
rect 3050 1334 3062 1336
rect 3018 1016 3020 1024
rect 3028 1016 3030 1024
rect 3018 1014 3030 1016
rect 2912 1006 2916 1014
rect 2924 1006 2928 1014
rect 2936 1006 2940 1014
rect 2948 1006 2952 1014
rect 2960 1006 2964 1014
rect 2972 1006 2976 1014
rect 2570 476 2572 484
rect 2580 476 2582 484
rect 2570 474 2582 476
rect 2912 614 2976 1006
rect 3114 964 3126 2096
rect 3242 2124 3254 2126
rect 3242 2116 3244 2124
rect 3252 2116 3254 2124
rect 3114 956 3116 964
rect 3124 956 3126 964
rect 3114 954 3126 956
rect 3178 1444 3190 1446
rect 3178 1436 3180 1444
rect 3188 1436 3190 1444
rect 2912 606 2916 614
rect 2924 606 2928 614
rect 2936 606 2940 614
rect 2948 606 2952 614
rect 2960 606 2964 614
rect 2972 606 2976 614
rect 1408 406 1412 414
rect 1420 406 1424 414
rect 1432 406 1436 414
rect 1444 406 1448 414
rect 1456 406 1460 414
rect 1468 406 1472 414
rect 1034 176 1036 184
rect 1044 176 1046 184
rect 1034 174 1046 176
rect 810 156 812 164
rect 820 156 822 164
rect 810 154 822 156
rect 1408 14 1472 406
rect 1866 344 1878 346
rect 1866 336 1868 344
rect 1876 336 1878 344
rect 1866 326 1878 336
rect 1834 314 1878 326
rect 1962 344 1974 346
rect 1962 336 1964 344
rect 1972 336 1974 344
rect 1834 284 1846 314
rect 1834 276 1836 284
rect 1844 276 1846 284
rect 1834 274 1846 276
rect 1962 284 1974 336
rect 1962 276 1964 284
rect 1972 276 1974 284
rect 1962 274 1974 276
rect 2090 324 2102 326
rect 2090 316 2092 324
rect 2100 316 2102 324
rect 2090 264 2102 316
rect 2090 256 2092 264
rect 2100 256 2102 264
rect 2090 254 2102 256
rect 2282 324 2294 326
rect 2282 316 2284 324
rect 2292 316 2294 324
rect 2282 184 2294 316
rect 2282 176 2284 184
rect 2292 176 2294 184
rect 2282 174 2294 176
rect 2912 214 2976 606
rect 3178 244 3190 1436
rect 3242 1284 3254 2116
rect 3370 2044 3382 2876
rect 3370 2036 3372 2044
rect 3380 2036 3382 2044
rect 3370 2034 3382 2036
rect 3402 2844 3414 2846
rect 3402 2836 3404 2844
rect 3412 2836 3414 2844
rect 3370 1864 3382 1866
rect 3370 1856 3372 1864
rect 3380 1856 3382 1864
rect 3370 1764 3382 1856
rect 3370 1756 3372 1764
rect 3380 1756 3382 1764
rect 3370 1504 3382 1756
rect 3402 1744 3414 2836
rect 3434 2624 3446 2626
rect 3434 2616 3436 2624
rect 3444 2616 3446 2624
rect 3434 1784 3446 2616
rect 3466 2364 3478 2896
rect 3466 2356 3468 2364
rect 3476 2356 3478 2364
rect 3466 2354 3478 2356
rect 3530 2304 3542 4496
rect 3594 3984 3606 4696
rect 3594 3976 3596 3984
rect 3604 3976 3606 3984
rect 3594 3974 3606 3976
rect 3626 4124 3638 4796
rect 3786 4584 3798 4956
rect 4010 4624 4022 5296
rect 4416 5214 4480 5416
rect 5920 5414 5984 5416
rect 5920 5406 5924 5414
rect 5932 5406 5936 5414
rect 5944 5406 5948 5414
rect 5956 5406 5960 5414
rect 5968 5406 5972 5414
rect 5980 5406 5984 5414
rect 5642 5404 5654 5406
rect 5642 5396 5644 5404
rect 5652 5396 5654 5404
rect 5322 5364 5398 5366
rect 5322 5356 5324 5364
rect 5332 5356 5398 5364
rect 5322 5354 5398 5356
rect 4416 5206 4420 5214
rect 4428 5206 4432 5214
rect 4440 5206 4444 5214
rect 4452 5206 4456 5214
rect 4464 5206 4468 5214
rect 4476 5206 4480 5214
rect 4010 4616 4012 4624
rect 4020 4616 4022 4624
rect 4010 4614 4022 4616
rect 4042 4944 4054 4946
rect 4042 4936 4044 4944
rect 4052 4936 4054 4944
rect 3786 4576 3788 4584
rect 3796 4576 3798 4584
rect 3786 4574 3798 4576
rect 3946 4424 3958 4426
rect 3946 4416 3948 4424
rect 3956 4416 3958 4424
rect 3626 4116 3628 4124
rect 3636 4116 3638 4124
rect 3594 3804 3606 3806
rect 3594 3796 3596 3804
rect 3604 3796 3606 3804
rect 3594 3644 3606 3796
rect 3594 3636 3596 3644
rect 3604 3636 3606 3644
rect 3594 3634 3606 3636
rect 3594 3304 3606 3306
rect 3594 3296 3596 3304
rect 3604 3296 3606 3304
rect 3594 3264 3606 3296
rect 3594 3256 3596 3264
rect 3604 3256 3606 3264
rect 3594 3254 3606 3256
rect 3530 2296 3532 2304
rect 3540 2296 3542 2304
rect 3530 2294 3542 2296
rect 3562 2304 3574 2306
rect 3562 2296 3564 2304
rect 3572 2296 3574 2304
rect 3530 2264 3542 2266
rect 3530 2256 3532 2264
rect 3540 2256 3542 2264
rect 3434 1776 3436 1784
rect 3444 1776 3446 1784
rect 3434 1774 3446 1776
rect 3498 1844 3510 1846
rect 3498 1836 3500 1844
rect 3508 1836 3510 1844
rect 3402 1736 3404 1744
rect 3412 1736 3414 1744
rect 3402 1734 3414 1736
rect 3370 1496 3372 1504
rect 3380 1496 3382 1504
rect 3370 1494 3382 1496
rect 3434 1504 3446 1506
rect 3434 1496 3436 1504
rect 3444 1496 3446 1504
rect 3242 1276 3244 1284
rect 3252 1276 3254 1284
rect 3242 1274 3254 1276
rect 3338 1344 3350 1346
rect 3338 1336 3340 1344
rect 3348 1336 3350 1344
rect 3210 1264 3222 1266
rect 3210 1256 3212 1264
rect 3220 1256 3222 1264
rect 3210 324 3222 1256
rect 3210 316 3212 324
rect 3220 316 3222 324
rect 3210 314 3222 316
rect 3338 264 3350 1336
rect 3434 1264 3446 1496
rect 3434 1256 3436 1264
rect 3444 1256 3446 1264
rect 3434 1254 3446 1256
rect 3498 1204 3510 1836
rect 3530 1784 3542 2256
rect 3530 1776 3532 1784
rect 3540 1776 3542 1784
rect 3530 1774 3542 1776
rect 3498 1196 3500 1204
rect 3508 1196 3510 1204
rect 3498 1194 3510 1196
rect 3530 1744 3542 1746
rect 3530 1736 3532 1744
rect 3540 1736 3542 1744
rect 3466 1124 3478 1126
rect 3466 1116 3468 1124
rect 3476 1116 3478 1124
rect 3370 984 3382 986
rect 3370 976 3372 984
rect 3380 976 3382 984
rect 3370 944 3382 976
rect 3370 936 3372 944
rect 3380 936 3382 944
rect 3370 934 3382 936
rect 3338 256 3340 264
rect 3348 256 3350 264
rect 3338 254 3350 256
rect 3178 236 3180 244
rect 3188 236 3190 244
rect 3178 234 3190 236
rect 2912 206 2916 214
rect 2924 206 2928 214
rect 2936 206 2940 214
rect 2948 206 2952 214
rect 2960 206 2964 214
rect 2972 206 2976 214
rect 1408 6 1412 14
rect 1420 6 1424 14
rect 1432 6 1436 14
rect 1444 6 1448 14
rect 1456 6 1460 14
rect 1468 6 1472 14
rect 1408 -10 1472 6
rect 2912 -10 2976 206
rect 3466 24 3478 1116
rect 3530 1084 3542 1736
rect 3562 1684 3574 2296
rect 3626 2124 3638 4116
rect 3722 4264 3734 4266
rect 3722 4256 3724 4264
rect 3732 4256 3734 4264
rect 3690 3764 3702 3766
rect 3690 3756 3692 3764
rect 3700 3756 3702 3764
rect 3690 3364 3702 3756
rect 3722 3624 3734 4256
rect 3882 4124 3894 4126
rect 3882 4116 3884 4124
rect 3892 4116 3894 4124
rect 3882 3884 3894 4116
rect 3882 3876 3884 3884
rect 3892 3876 3894 3884
rect 3850 3784 3862 3786
rect 3850 3776 3852 3784
rect 3860 3776 3862 3784
rect 3850 3724 3862 3776
rect 3850 3716 3852 3724
rect 3860 3716 3862 3724
rect 3850 3714 3862 3716
rect 3722 3616 3724 3624
rect 3732 3616 3734 3624
rect 3722 3614 3734 3616
rect 3850 3524 3862 3526
rect 3850 3516 3852 3524
rect 3860 3516 3862 3524
rect 3690 3356 3692 3364
rect 3700 3356 3702 3364
rect 3690 3354 3702 3356
rect 3722 3364 3734 3366
rect 3722 3356 3724 3364
rect 3732 3356 3734 3364
rect 3658 3264 3670 3266
rect 3658 3256 3660 3264
rect 3668 3256 3670 3264
rect 3658 2244 3670 3256
rect 3722 2984 3734 3356
rect 3722 2976 3724 2984
rect 3732 2976 3734 2984
rect 3722 2974 3734 2976
rect 3818 2904 3830 2906
rect 3818 2896 3820 2904
rect 3828 2896 3830 2904
rect 3754 2784 3766 2786
rect 3754 2776 3756 2784
rect 3764 2776 3766 2784
rect 3722 2764 3734 2766
rect 3722 2756 3724 2764
rect 3732 2756 3734 2764
rect 3690 2724 3702 2726
rect 3690 2716 3692 2724
rect 3700 2716 3702 2724
rect 3690 2484 3702 2716
rect 3722 2724 3734 2756
rect 3722 2716 3724 2724
rect 3732 2716 3734 2724
rect 3722 2714 3734 2716
rect 3690 2476 3692 2484
rect 3700 2476 3702 2484
rect 3690 2284 3702 2476
rect 3690 2276 3692 2284
rect 3700 2276 3702 2284
rect 3690 2274 3702 2276
rect 3722 2664 3734 2666
rect 3722 2656 3724 2664
rect 3732 2656 3734 2664
rect 3658 2236 3660 2244
rect 3668 2236 3670 2244
rect 3658 2234 3670 2236
rect 3690 2244 3702 2246
rect 3690 2236 3692 2244
rect 3700 2236 3702 2244
rect 3690 2204 3702 2236
rect 3690 2196 3692 2204
rect 3700 2196 3702 2204
rect 3690 2194 3702 2196
rect 3626 2116 3628 2124
rect 3636 2116 3638 2124
rect 3562 1676 3564 1684
rect 3572 1676 3574 1684
rect 3562 1674 3574 1676
rect 3594 2044 3606 2046
rect 3594 2036 3596 2044
rect 3604 2036 3606 2044
rect 3594 1244 3606 2036
rect 3626 1504 3638 2116
rect 3722 2124 3734 2656
rect 3754 2244 3766 2776
rect 3786 2744 3798 2746
rect 3786 2736 3788 2744
rect 3796 2736 3798 2744
rect 3786 2564 3798 2736
rect 3786 2556 3788 2564
rect 3796 2556 3798 2564
rect 3786 2554 3798 2556
rect 3818 2524 3830 2896
rect 3850 2904 3862 3516
rect 3850 2896 3852 2904
rect 3860 2896 3862 2904
rect 3850 2894 3862 2896
rect 3882 3484 3894 3876
rect 3946 3544 3958 4416
rect 3946 3536 3948 3544
rect 3956 3536 3958 3544
rect 3946 3534 3958 3536
rect 3882 3476 3884 3484
rect 3892 3476 3894 3484
rect 3882 2964 3894 3476
rect 3882 2956 3884 2964
rect 3892 2956 3894 2964
rect 3818 2516 3820 2524
rect 3828 2516 3830 2524
rect 3818 2514 3830 2516
rect 3850 2664 3862 2666
rect 3850 2656 3852 2664
rect 3860 2656 3862 2664
rect 3754 2236 3756 2244
rect 3764 2236 3766 2244
rect 3754 2234 3766 2236
rect 3850 2144 3862 2656
rect 3882 2364 3894 2956
rect 4010 2984 4022 2986
rect 4010 2976 4012 2984
rect 4020 2976 4022 2984
rect 3914 2684 3926 2686
rect 3914 2676 3916 2684
rect 3924 2676 3926 2684
rect 3914 2544 3926 2676
rect 4010 2664 4022 2976
rect 4010 2656 4012 2664
rect 4020 2656 4022 2664
rect 4010 2654 4022 2656
rect 3914 2536 3916 2544
rect 3924 2536 3926 2544
rect 3914 2534 3926 2536
rect 3978 2604 3990 2606
rect 3978 2596 3980 2604
rect 3988 2596 3990 2604
rect 3882 2356 3884 2364
rect 3892 2356 3894 2364
rect 3882 2354 3894 2356
rect 3914 2404 3926 2406
rect 3914 2396 3916 2404
rect 3924 2396 3926 2404
rect 3914 2244 3926 2396
rect 3914 2236 3916 2244
rect 3924 2236 3926 2244
rect 3914 2234 3926 2236
rect 3946 2264 3958 2266
rect 3946 2256 3948 2264
rect 3956 2256 3958 2264
rect 3850 2136 3852 2144
rect 3860 2136 3862 2144
rect 3850 2134 3862 2136
rect 3722 2116 3724 2124
rect 3732 2116 3734 2124
rect 3722 2114 3734 2116
rect 3786 2124 3798 2126
rect 3786 2116 3788 2124
rect 3796 2116 3798 2124
rect 3786 2024 3798 2116
rect 3786 2016 3788 2024
rect 3796 2016 3798 2024
rect 3786 2014 3798 2016
rect 3722 1964 3734 1966
rect 3722 1956 3724 1964
rect 3732 1956 3734 1964
rect 3722 1924 3734 1956
rect 3722 1916 3724 1924
rect 3732 1916 3734 1924
rect 3722 1914 3734 1916
rect 3722 1884 3734 1886
rect 3722 1876 3724 1884
rect 3732 1876 3734 1884
rect 3690 1864 3702 1866
rect 3690 1856 3692 1864
rect 3700 1856 3702 1864
rect 3690 1684 3702 1856
rect 3690 1676 3692 1684
rect 3700 1676 3702 1684
rect 3690 1674 3702 1676
rect 3626 1496 3628 1504
rect 3636 1496 3638 1504
rect 3626 1404 3638 1496
rect 3722 1504 3734 1876
rect 3914 1764 3926 1766
rect 3914 1756 3916 1764
rect 3924 1756 3926 1764
rect 3786 1724 3798 1726
rect 3786 1716 3788 1724
rect 3796 1716 3798 1724
rect 3786 1684 3798 1716
rect 3786 1676 3788 1684
rect 3796 1676 3798 1684
rect 3786 1674 3798 1676
rect 3722 1496 3724 1504
rect 3732 1496 3734 1504
rect 3722 1494 3734 1496
rect 3786 1644 3798 1646
rect 3786 1636 3788 1644
rect 3796 1636 3798 1644
rect 3626 1396 3628 1404
rect 3636 1396 3638 1404
rect 3626 1394 3638 1396
rect 3786 1344 3798 1636
rect 3914 1584 3926 1756
rect 3914 1576 3916 1584
rect 3924 1576 3926 1584
rect 3914 1574 3926 1576
rect 3946 1584 3958 2256
rect 3978 1924 3990 2596
rect 4010 2404 4022 2406
rect 4010 2396 4012 2404
rect 4020 2396 4022 2404
rect 4010 2204 4022 2396
rect 4042 2364 4054 4936
rect 4416 4814 4480 5206
rect 5322 5324 5334 5326
rect 5322 5316 5324 5324
rect 5332 5316 5334 5324
rect 5194 5164 5206 5166
rect 5194 5156 5196 5164
rect 5204 5156 5206 5164
rect 4714 5144 4726 5146
rect 4714 5136 4716 5144
rect 4724 5136 4726 5144
rect 4650 5124 4662 5126
rect 4650 5116 4652 5124
rect 4660 5116 4662 5124
rect 4618 5004 4630 5006
rect 4618 4996 4620 5004
rect 4628 4996 4630 5004
rect 4618 4924 4630 4996
rect 4618 4916 4620 4924
rect 4628 4916 4630 4924
rect 4618 4914 4630 4916
rect 4416 4806 4420 4814
rect 4428 4806 4432 4814
rect 4440 4806 4444 4814
rect 4452 4806 4456 4814
rect 4464 4806 4468 4814
rect 4476 4806 4480 4814
rect 4106 4744 4118 4746
rect 4106 4736 4108 4744
rect 4116 4736 4118 4744
rect 4106 4364 4118 4736
rect 4106 4356 4108 4364
rect 4116 4356 4118 4364
rect 4106 4354 4118 4356
rect 4416 4414 4480 4806
rect 4522 4804 4534 4806
rect 4522 4796 4524 4804
rect 4532 4796 4534 4804
rect 4522 4764 4534 4796
rect 4522 4756 4524 4764
rect 4532 4756 4534 4764
rect 4522 4754 4534 4756
rect 4522 4644 4534 4646
rect 4522 4636 4524 4644
rect 4532 4636 4534 4644
rect 4522 4424 4534 4636
rect 4650 4584 4662 5116
rect 4650 4576 4652 4584
rect 4660 4576 4662 4584
rect 4650 4574 4662 4576
rect 4682 4684 4694 4686
rect 4682 4676 4684 4684
rect 4692 4676 4694 4684
rect 4522 4416 4524 4424
rect 4532 4416 4534 4424
rect 4522 4414 4534 4416
rect 4586 4524 4598 4526
rect 4586 4516 4588 4524
rect 4596 4516 4598 4524
rect 4586 4444 4598 4516
rect 4586 4436 4588 4444
rect 4596 4436 4598 4444
rect 4416 4406 4420 4414
rect 4428 4406 4432 4414
rect 4440 4406 4444 4414
rect 4452 4406 4456 4414
rect 4464 4406 4468 4414
rect 4476 4406 4480 4414
rect 4362 4144 4374 4146
rect 4362 4136 4364 4144
rect 4372 4136 4374 4144
rect 4106 3924 4118 3926
rect 4106 3916 4108 3924
rect 4116 3916 4118 3924
rect 4106 3524 4118 3916
rect 4106 3516 4108 3524
rect 4116 3516 4118 3524
rect 4106 3514 4118 3516
rect 4202 3804 4214 3806
rect 4202 3796 4204 3804
rect 4212 3796 4214 3804
rect 4074 3304 4086 3306
rect 4074 3296 4076 3304
rect 4084 3296 4086 3304
rect 4074 2884 4086 3296
rect 4074 2876 4076 2884
rect 4084 2876 4086 2884
rect 4074 2874 4086 2876
rect 4138 3204 4150 3206
rect 4138 3196 4140 3204
rect 4148 3196 4150 3204
rect 4074 2744 4086 2746
rect 4074 2736 4076 2744
rect 4084 2736 4086 2744
rect 4074 2504 4086 2736
rect 4138 2704 4150 3196
rect 4202 3144 4214 3796
rect 4298 3804 4310 3806
rect 4298 3796 4300 3804
rect 4308 3796 4310 3804
rect 4266 3764 4278 3766
rect 4266 3756 4268 3764
rect 4276 3756 4278 3764
rect 4266 3724 4278 3756
rect 4266 3716 4268 3724
rect 4276 3716 4278 3724
rect 4266 3714 4278 3716
rect 4298 3504 4310 3796
rect 4298 3496 4300 3504
rect 4308 3496 4310 3504
rect 4298 3494 4310 3496
rect 4202 3136 4204 3144
rect 4212 3136 4214 3144
rect 4202 3104 4214 3136
rect 4202 3096 4204 3104
rect 4212 3096 4214 3104
rect 4138 2696 4140 2704
rect 4148 2696 4150 2704
rect 4138 2694 4150 2696
rect 4170 3084 4182 3086
rect 4170 3076 4172 3084
rect 4180 3076 4182 3084
rect 4170 2924 4182 3076
rect 4202 3064 4214 3096
rect 4202 3056 4204 3064
rect 4212 3056 4214 3064
rect 4202 3054 4214 3056
rect 4234 3324 4246 3326
rect 4234 3316 4236 3324
rect 4244 3316 4246 3324
rect 4170 2916 4172 2924
rect 4180 2916 4182 2924
rect 4138 2664 4150 2666
rect 4138 2656 4140 2664
rect 4148 2656 4150 2664
rect 4138 2646 4150 2656
rect 4106 2634 4150 2646
rect 4106 2604 4118 2634
rect 4106 2596 4108 2604
rect 4116 2596 4118 2604
rect 4106 2594 4118 2596
rect 4138 2604 4150 2606
rect 4138 2596 4140 2604
rect 4148 2596 4150 2604
rect 4074 2496 4076 2504
rect 4084 2496 4086 2504
rect 4074 2494 4086 2496
rect 4106 2564 4118 2566
rect 4106 2556 4108 2564
rect 4116 2556 4118 2564
rect 4106 2464 4118 2556
rect 4106 2456 4108 2464
rect 4116 2456 4118 2464
rect 4106 2454 4118 2456
rect 4138 2464 4150 2596
rect 4138 2456 4140 2464
rect 4148 2456 4150 2464
rect 4138 2454 4150 2456
rect 4042 2356 4044 2364
rect 4052 2356 4054 2364
rect 4042 2354 4054 2356
rect 4074 2364 4086 2366
rect 4074 2356 4076 2364
rect 4084 2356 4086 2364
rect 4074 2244 4086 2356
rect 4074 2236 4076 2244
rect 4084 2236 4086 2244
rect 4074 2234 4086 2236
rect 4010 2196 4012 2204
rect 4020 2196 4022 2204
rect 4010 2194 4022 2196
rect 4074 2164 4086 2166
rect 4074 2156 4076 2164
rect 4084 2156 4086 2164
rect 3978 1916 3980 1924
rect 3988 1916 3990 1924
rect 3978 1914 3990 1916
rect 4010 2124 4022 2126
rect 4010 2116 4012 2124
rect 4020 2116 4022 2124
rect 4010 1764 4022 2116
rect 4074 2084 4086 2156
rect 4074 2076 4076 2084
rect 4084 2076 4086 2084
rect 4074 2074 4086 2076
rect 4138 2164 4150 2166
rect 4138 2156 4140 2164
rect 4148 2156 4150 2164
rect 4138 1924 4150 2156
rect 4138 1916 4140 1924
rect 4148 1916 4150 1924
rect 4138 1914 4150 1916
rect 4010 1756 4012 1764
rect 4020 1756 4022 1764
rect 4010 1754 4022 1756
rect 4074 1864 4086 1866
rect 4074 1856 4076 1864
rect 4084 1856 4086 1864
rect 4074 1664 4086 1856
rect 4138 1864 4150 1866
rect 4138 1856 4140 1864
rect 4148 1856 4150 1864
rect 4138 1724 4150 1856
rect 4138 1716 4140 1724
rect 4148 1716 4150 1724
rect 4138 1714 4150 1716
rect 4074 1656 4076 1664
rect 4084 1656 4086 1664
rect 4074 1654 4086 1656
rect 4138 1624 4150 1626
rect 4138 1616 4140 1624
rect 4148 1616 4150 1624
rect 3946 1576 3948 1584
rect 3956 1576 3958 1584
rect 3946 1574 3958 1576
rect 3978 1584 3990 1586
rect 3978 1576 3980 1584
rect 3988 1576 3990 1584
rect 3978 1544 3990 1576
rect 4138 1564 4150 1616
rect 4138 1556 4140 1564
rect 4148 1556 4150 1564
rect 4138 1554 4150 1556
rect 3978 1536 3980 1544
rect 3988 1536 3990 1544
rect 3978 1534 3990 1536
rect 3818 1524 3830 1526
rect 3818 1516 3820 1524
rect 3828 1516 3830 1524
rect 3818 1404 3830 1516
rect 3818 1396 3820 1404
rect 3828 1396 3830 1404
rect 3818 1394 3830 1396
rect 4074 1444 4086 1446
rect 4074 1436 4076 1444
rect 4084 1436 4086 1444
rect 3786 1336 3788 1344
rect 3796 1336 3798 1344
rect 3786 1334 3798 1336
rect 3594 1236 3596 1244
rect 3604 1236 3606 1244
rect 3594 1234 3606 1236
rect 3946 1224 3958 1226
rect 3946 1216 3948 1224
rect 3956 1216 3958 1224
rect 3946 1164 3958 1216
rect 3946 1156 3948 1164
rect 3956 1156 3958 1164
rect 3946 1154 3958 1156
rect 3530 1076 3532 1084
rect 3540 1076 3542 1084
rect 3530 1074 3542 1076
rect 4074 1064 4086 1436
rect 4170 1164 4182 2916
rect 4202 3004 4214 3006
rect 4202 2996 4204 3004
rect 4212 2996 4214 3004
rect 4202 2904 4214 2996
rect 4202 2896 4204 2904
rect 4212 2896 4214 2904
rect 4202 2894 4214 2896
rect 4202 2704 4214 2706
rect 4202 2696 4204 2704
rect 4212 2696 4214 2704
rect 4202 1884 4214 2696
rect 4202 1876 4204 1884
rect 4212 1876 4214 1884
rect 4202 1874 4214 1876
rect 4234 2544 4246 3316
rect 4266 3304 4278 3306
rect 4266 3296 4268 3304
rect 4276 3296 4278 3304
rect 4266 2804 4278 3296
rect 4330 3064 4342 3066
rect 4330 3056 4332 3064
rect 4340 3056 4342 3064
rect 4266 2796 4268 2804
rect 4276 2796 4278 2804
rect 4266 2794 4278 2796
rect 4298 3024 4310 3026
rect 4298 3016 4300 3024
rect 4308 3016 4310 3024
rect 4298 2744 4310 3016
rect 4298 2736 4300 2744
rect 4308 2736 4310 2744
rect 4298 2734 4310 2736
rect 4330 2944 4342 3056
rect 4362 3004 4374 4136
rect 4362 2996 4364 3004
rect 4372 2996 4374 3004
rect 4362 2994 4374 2996
rect 4416 4014 4480 4406
rect 4416 4006 4420 4014
rect 4428 4006 4432 4014
rect 4440 4006 4444 4014
rect 4452 4006 4456 4014
rect 4464 4006 4468 4014
rect 4476 4006 4480 4014
rect 4416 3614 4480 4006
rect 4586 3984 4598 4436
rect 4682 4164 4694 4676
rect 4714 4684 4726 5136
rect 5162 5084 5174 5086
rect 5162 5076 5164 5084
rect 5172 5076 5174 5084
rect 5098 4964 5110 4966
rect 5098 4956 5100 4964
rect 5108 4956 5110 4964
rect 4874 4924 4886 4926
rect 4874 4916 4876 4924
rect 4884 4916 4886 4924
rect 4714 4676 4716 4684
rect 4724 4676 4726 4684
rect 4714 4674 4726 4676
rect 4778 4764 4790 4766
rect 4778 4756 4780 4764
rect 4788 4756 4790 4764
rect 4778 4604 4790 4756
rect 4778 4596 4780 4604
rect 4788 4596 4790 4604
rect 4778 4594 4790 4596
rect 4874 4584 4886 4916
rect 5098 4904 5110 4956
rect 5098 4896 5100 4904
rect 5108 4896 5110 4904
rect 5098 4894 5110 4896
rect 5002 4864 5014 4866
rect 5002 4856 5004 4864
rect 5012 4856 5014 4864
rect 4874 4576 4876 4584
rect 4884 4576 4886 4584
rect 4874 4574 4886 4576
rect 4938 4704 4950 4706
rect 4938 4696 4940 4704
rect 4948 4696 4950 4704
rect 4682 4156 4684 4164
rect 4692 4156 4694 4164
rect 4682 4154 4694 4156
rect 4874 4284 4886 4286
rect 4874 4276 4876 4284
rect 4884 4276 4886 4284
rect 4586 3976 4588 3984
rect 4596 3976 4598 3984
rect 4586 3974 4598 3976
rect 4416 3606 4420 3614
rect 4428 3606 4432 3614
rect 4440 3606 4444 3614
rect 4452 3606 4456 3614
rect 4464 3606 4468 3614
rect 4476 3606 4480 3614
rect 4416 3214 4480 3606
rect 4416 3206 4420 3214
rect 4428 3206 4432 3214
rect 4440 3206 4444 3214
rect 4452 3206 4456 3214
rect 4464 3206 4468 3214
rect 4476 3206 4480 3214
rect 4330 2936 4332 2944
rect 4340 2936 4342 2944
rect 4266 2684 4278 2686
rect 4266 2676 4268 2684
rect 4276 2676 4278 2684
rect 4266 2624 4278 2676
rect 4266 2616 4268 2624
rect 4276 2616 4278 2624
rect 4266 2614 4278 2616
rect 4234 2536 4236 2544
rect 4244 2536 4246 2544
rect 4234 1904 4246 2536
rect 4266 2504 4278 2506
rect 4266 2496 4268 2504
rect 4276 2496 4278 2504
rect 4266 2184 4278 2496
rect 4298 2484 4310 2486
rect 4298 2476 4300 2484
rect 4308 2476 4310 2484
rect 4298 2424 4310 2476
rect 4298 2416 4300 2424
rect 4308 2416 4310 2424
rect 4298 2414 4310 2416
rect 4266 2176 4268 2184
rect 4276 2176 4278 2184
rect 4266 2174 4278 2176
rect 4298 2224 4310 2226
rect 4298 2216 4300 2224
rect 4308 2216 4310 2224
rect 4234 1896 4236 1904
rect 4244 1896 4246 1904
rect 4202 1724 4214 1726
rect 4202 1716 4204 1724
rect 4212 1716 4214 1724
rect 4202 1604 4214 1716
rect 4202 1596 4204 1604
rect 4212 1596 4214 1604
rect 4202 1594 4214 1596
rect 4234 1384 4246 1896
rect 4266 2124 4278 2126
rect 4266 2116 4268 2124
rect 4276 2116 4278 2124
rect 4266 1864 4278 2116
rect 4298 2104 4310 2216
rect 4298 2096 4300 2104
rect 4308 2096 4310 2104
rect 4298 2094 4310 2096
rect 4266 1856 4268 1864
rect 4276 1856 4278 1864
rect 4266 1854 4278 1856
rect 4298 1884 4310 1886
rect 4298 1876 4300 1884
rect 4308 1876 4310 1884
rect 4298 1824 4310 1876
rect 4298 1816 4300 1824
rect 4308 1816 4310 1824
rect 4298 1814 4310 1816
rect 4298 1784 4310 1786
rect 4298 1776 4300 1784
rect 4308 1776 4310 1784
rect 4298 1484 4310 1776
rect 4298 1476 4300 1484
rect 4308 1476 4310 1484
rect 4298 1474 4310 1476
rect 4234 1376 4236 1384
rect 4244 1376 4246 1384
rect 4234 1374 4246 1376
rect 4298 1424 4310 1426
rect 4298 1416 4300 1424
rect 4308 1416 4310 1424
rect 4170 1156 4172 1164
rect 4180 1156 4182 1164
rect 4170 1154 4182 1156
rect 4074 1056 4076 1064
rect 4084 1056 4086 1064
rect 4074 1054 4086 1056
rect 4106 1124 4118 1126
rect 4106 1116 4108 1124
rect 4116 1116 4118 1124
rect 4042 1024 4054 1026
rect 4042 1016 4044 1024
rect 4052 1016 4054 1024
rect 3658 1004 3670 1006
rect 3658 996 3660 1004
rect 3668 996 3670 1004
rect 3466 16 3468 24
rect 3476 16 3478 24
rect 3466 14 3478 16
rect 3594 544 3606 546
rect 3594 536 3596 544
rect 3604 536 3606 544
rect 3594 24 3606 536
rect 3594 16 3596 24
rect 3604 16 3606 24
rect 3594 14 3606 16
rect 3658 24 3670 996
rect 3978 824 3990 826
rect 3978 816 3980 824
rect 3988 816 3990 824
rect 3946 724 3958 726
rect 3946 716 3948 724
rect 3956 716 3958 724
rect 3850 704 3862 706
rect 3850 696 3852 704
rect 3860 696 3862 704
rect 3754 644 3766 646
rect 3754 636 3756 644
rect 3764 636 3766 644
rect 3754 104 3766 636
rect 3850 384 3862 696
rect 3946 544 3958 716
rect 3946 536 3948 544
rect 3956 536 3958 544
rect 3946 534 3958 536
rect 3978 544 3990 816
rect 4042 764 4054 1016
rect 4042 756 4044 764
rect 4052 756 4054 764
rect 4042 754 4054 756
rect 3978 536 3980 544
rect 3988 536 3990 544
rect 3978 534 3990 536
rect 4042 664 4054 666
rect 4042 656 4044 664
rect 4052 656 4054 664
rect 3850 376 3852 384
rect 3860 376 3862 384
rect 3850 374 3862 376
rect 3882 344 3894 346
rect 3882 336 3884 344
rect 3892 336 3894 344
rect 3882 184 3894 336
rect 4042 284 4054 656
rect 4106 624 4118 1116
rect 4202 1104 4214 1106
rect 4202 1096 4204 1104
rect 4212 1096 4214 1104
rect 4106 616 4108 624
rect 4116 616 4118 624
rect 4106 614 4118 616
rect 4170 1084 4182 1086
rect 4170 1076 4172 1084
rect 4180 1076 4182 1084
rect 4170 484 4182 1076
rect 4202 644 4214 1096
rect 4234 784 4246 786
rect 4234 776 4236 784
rect 4244 776 4246 784
rect 4234 684 4246 776
rect 4234 676 4236 684
rect 4244 676 4246 684
rect 4234 674 4246 676
rect 4202 636 4204 644
rect 4212 636 4214 644
rect 4202 634 4214 636
rect 4170 476 4172 484
rect 4180 476 4182 484
rect 4170 474 4182 476
rect 4298 364 4310 1416
rect 4330 744 4342 2936
rect 4416 2814 4480 3206
rect 4554 3704 4566 3706
rect 4554 3696 4556 3704
rect 4564 3696 4566 3704
rect 4554 2964 4566 3696
rect 4618 3504 4630 3506
rect 4618 3496 4620 3504
rect 4628 3496 4630 3504
rect 4554 2956 4556 2964
rect 4564 2956 4566 2964
rect 4554 2954 4566 2956
rect 4586 3164 4598 3166
rect 4586 3156 4588 3164
rect 4596 3156 4598 3164
rect 4416 2806 4420 2814
rect 4428 2806 4432 2814
rect 4440 2806 4444 2814
rect 4452 2806 4456 2814
rect 4464 2806 4468 2814
rect 4476 2806 4480 2814
rect 4362 2464 4374 2466
rect 4362 2456 4364 2464
rect 4372 2456 4374 2464
rect 4362 2144 4374 2456
rect 4362 2136 4364 2144
rect 4372 2136 4374 2144
rect 4362 2134 4374 2136
rect 4416 2414 4480 2806
rect 4416 2406 4420 2414
rect 4428 2406 4432 2414
rect 4440 2406 4444 2414
rect 4452 2406 4456 2414
rect 4464 2406 4468 2414
rect 4476 2406 4480 2414
rect 4416 2014 4480 2406
rect 4522 2804 4534 2806
rect 4522 2796 4524 2804
rect 4532 2796 4534 2804
rect 4522 2184 4534 2796
rect 4586 2664 4598 3156
rect 4618 2864 4630 3496
rect 4618 2856 4620 2864
rect 4628 2856 4630 2864
rect 4618 2854 4630 2856
rect 4714 3104 4726 3106
rect 4714 3096 4716 3104
rect 4724 3096 4726 3104
rect 4714 2904 4726 3096
rect 4874 2924 4886 4276
rect 4906 3824 4918 3826
rect 4906 3816 4908 3824
rect 4916 3816 4918 3824
rect 4906 3684 4918 3816
rect 4938 3724 4950 4696
rect 5002 4444 5014 4856
rect 5162 4784 5174 5076
rect 5162 4776 5164 4784
rect 5172 4776 5174 4784
rect 5002 4436 5004 4444
rect 5012 4436 5014 4444
rect 5002 4434 5014 4436
rect 5034 4684 5046 4686
rect 5034 4676 5036 4684
rect 5044 4676 5046 4684
rect 4938 3716 4940 3724
rect 4948 3716 4950 3724
rect 4938 3714 4950 3716
rect 5034 3724 5046 4676
rect 5162 4524 5174 4776
rect 5194 4724 5206 5156
rect 5322 5024 5334 5316
rect 5386 5324 5398 5354
rect 5386 5316 5388 5324
rect 5396 5316 5398 5324
rect 5386 5314 5398 5316
rect 5418 5364 5430 5366
rect 5418 5356 5420 5364
rect 5428 5356 5430 5364
rect 5322 5016 5324 5024
rect 5332 5016 5334 5024
rect 5322 5014 5334 5016
rect 5354 5304 5366 5306
rect 5354 5296 5356 5304
rect 5364 5296 5366 5304
rect 5194 4716 5196 4724
rect 5204 4716 5206 4724
rect 5194 4714 5206 4716
rect 5258 4924 5270 4926
rect 5258 4916 5260 4924
rect 5268 4916 5270 4924
rect 5162 4516 5164 4524
rect 5172 4516 5174 4524
rect 5162 4514 5174 4516
rect 5258 4484 5270 4916
rect 5354 4844 5366 5296
rect 5418 5304 5430 5356
rect 5418 5296 5420 5304
rect 5428 5296 5430 5304
rect 5418 5294 5430 5296
rect 5546 5104 5558 5106
rect 5546 5096 5548 5104
rect 5556 5096 5558 5104
rect 5482 5084 5494 5086
rect 5482 5076 5484 5084
rect 5492 5076 5494 5084
rect 5354 4836 5356 4844
rect 5364 4836 5366 4844
rect 5354 4834 5366 4836
rect 5386 4944 5398 4946
rect 5386 4936 5388 4944
rect 5396 4936 5398 4944
rect 5386 4664 5398 4936
rect 5482 4784 5494 5076
rect 5482 4776 5484 4784
rect 5492 4776 5494 4784
rect 5482 4774 5494 4776
rect 5386 4656 5388 4664
rect 5396 4656 5398 4664
rect 5386 4654 5398 4656
rect 5514 4744 5526 4746
rect 5514 4736 5516 4744
rect 5524 4736 5526 4744
rect 5258 4476 5260 4484
rect 5268 4476 5270 4484
rect 5258 4474 5270 4476
rect 5354 4504 5366 4506
rect 5354 4496 5356 4504
rect 5364 4496 5366 4504
rect 5130 4344 5142 4346
rect 5130 4336 5132 4344
rect 5140 4336 5142 4344
rect 5130 4184 5142 4336
rect 5130 4176 5132 4184
rect 5140 4176 5142 4184
rect 5130 4174 5142 4176
rect 5322 4344 5334 4346
rect 5322 4336 5324 4344
rect 5332 4336 5334 4344
rect 5322 3884 5334 4336
rect 5354 4264 5366 4496
rect 5514 4464 5526 4736
rect 5514 4456 5516 4464
rect 5524 4456 5526 4464
rect 5514 4454 5526 4456
rect 5546 4724 5558 5096
rect 5642 4984 5654 5396
rect 5802 5264 5814 5266
rect 5802 5256 5804 5264
rect 5812 5256 5814 5264
rect 5738 5144 5750 5146
rect 5738 5136 5740 5144
rect 5748 5136 5750 5144
rect 5642 4976 5644 4984
rect 5652 4976 5654 4984
rect 5642 4974 5654 4976
rect 5706 5124 5718 5126
rect 5706 5116 5708 5124
rect 5716 5116 5718 5124
rect 5610 4944 5622 4946
rect 5610 4936 5612 4944
rect 5620 4936 5622 4944
rect 5610 4824 5622 4936
rect 5706 4924 5718 5116
rect 5738 5064 5750 5136
rect 5738 5056 5740 5064
rect 5748 5056 5750 5064
rect 5738 5054 5750 5056
rect 5706 4916 5708 4924
rect 5716 4916 5718 4924
rect 5706 4914 5718 4916
rect 5802 4844 5814 5256
rect 5802 4836 5804 4844
rect 5812 4836 5814 4844
rect 5802 4834 5814 4836
rect 5920 5014 5984 5406
rect 5920 5006 5924 5014
rect 5932 5006 5936 5014
rect 5944 5006 5948 5014
rect 5956 5006 5960 5014
rect 5968 5006 5972 5014
rect 5980 5006 5984 5014
rect 5610 4816 5612 4824
rect 5620 4816 5622 4824
rect 5610 4814 5622 4816
rect 5546 4716 5548 4724
rect 5556 4716 5558 4724
rect 5450 4424 5462 4426
rect 5450 4416 5452 4424
rect 5460 4416 5462 4424
rect 5354 4256 5356 4264
rect 5364 4256 5366 4264
rect 5354 4254 5366 4256
rect 5386 4344 5398 4346
rect 5386 4336 5388 4344
rect 5396 4336 5398 4344
rect 5386 4144 5398 4336
rect 5386 4136 5388 4144
rect 5396 4136 5398 4144
rect 5386 4134 5398 4136
rect 5450 4104 5462 4416
rect 5450 4096 5452 4104
rect 5460 4096 5462 4104
rect 5450 4094 5462 4096
rect 5546 4304 5558 4716
rect 5866 4704 5878 4706
rect 5866 4696 5868 4704
rect 5876 4696 5878 4704
rect 5802 4684 5814 4686
rect 5802 4676 5804 4684
rect 5812 4676 5814 4684
rect 5610 4524 5622 4526
rect 5610 4516 5612 4524
rect 5620 4516 5622 4524
rect 5610 4444 5622 4516
rect 5610 4436 5612 4444
rect 5620 4436 5622 4444
rect 5546 4296 5548 4304
rect 5556 4296 5558 4304
rect 5322 3876 5324 3884
rect 5332 3876 5334 3884
rect 5322 3764 5334 3876
rect 5322 3756 5324 3764
rect 5332 3756 5334 3764
rect 5322 3754 5334 3756
rect 5418 3864 5430 3866
rect 5418 3856 5420 3864
rect 5428 3856 5430 3864
rect 5034 3716 5036 3724
rect 5044 3716 5046 3724
rect 5034 3714 5046 3716
rect 5194 3744 5206 3746
rect 5194 3736 5196 3744
rect 5204 3736 5206 3744
rect 4906 3676 4908 3684
rect 4916 3676 4918 3684
rect 4906 3674 4918 3676
rect 5098 3704 5110 3706
rect 5098 3696 5100 3704
rect 5108 3696 5110 3704
rect 5098 3664 5110 3696
rect 5098 3656 5100 3664
rect 5108 3656 5110 3664
rect 5098 3364 5110 3656
rect 5098 3356 5100 3364
rect 5108 3356 5110 3364
rect 5098 3354 5110 3356
rect 5162 3464 5174 3466
rect 5162 3456 5164 3464
rect 5172 3456 5174 3464
rect 5162 3104 5174 3456
rect 5162 3096 5164 3104
rect 5172 3096 5174 3104
rect 5162 3094 5174 3096
rect 5194 3084 5206 3736
rect 5386 3744 5398 3746
rect 5386 3736 5388 3744
rect 5396 3736 5398 3744
rect 5386 3164 5398 3736
rect 5418 3744 5430 3856
rect 5418 3736 5420 3744
rect 5428 3736 5430 3744
rect 5418 3734 5430 3736
rect 5386 3156 5388 3164
rect 5396 3156 5398 3164
rect 5386 3154 5398 3156
rect 5450 3364 5462 3366
rect 5450 3356 5452 3364
rect 5460 3356 5462 3364
rect 5450 3244 5462 3356
rect 5450 3236 5452 3244
rect 5460 3236 5462 3244
rect 5450 3104 5462 3236
rect 5450 3096 5452 3104
rect 5460 3096 5462 3104
rect 5450 3094 5462 3096
rect 5194 3076 5196 3084
rect 5204 3076 5206 3084
rect 5194 3074 5206 3076
rect 4874 2916 4876 2924
rect 4884 2916 4886 2924
rect 4874 2914 4886 2916
rect 5546 2924 5558 4296
rect 5578 4304 5590 4306
rect 5578 4296 5580 4304
rect 5588 4296 5590 4304
rect 5578 4204 5590 4296
rect 5578 4196 5580 4204
rect 5588 4196 5590 4204
rect 5578 4194 5590 4196
rect 5610 3784 5622 4436
rect 5642 4304 5654 4306
rect 5642 4296 5644 4304
rect 5652 4296 5654 4304
rect 5642 4244 5654 4296
rect 5770 4304 5782 4306
rect 5770 4296 5772 4304
rect 5780 4296 5782 4304
rect 5642 4236 5644 4244
rect 5652 4236 5654 4244
rect 5642 4234 5654 4236
rect 5738 4264 5750 4266
rect 5738 4256 5740 4264
rect 5748 4256 5750 4264
rect 5738 4204 5750 4256
rect 5738 4196 5740 4204
rect 5748 4196 5750 4204
rect 5610 3776 5612 3784
rect 5620 3776 5622 3784
rect 5610 3774 5622 3776
rect 5642 4144 5654 4146
rect 5642 4136 5644 4144
rect 5652 4136 5654 4144
rect 5546 2916 5548 2924
rect 5556 2916 5558 2924
rect 5546 2914 5558 2916
rect 5578 2924 5590 2926
rect 5578 2916 5580 2924
rect 5588 2916 5590 2924
rect 4714 2896 4716 2904
rect 4724 2896 4726 2904
rect 4586 2656 4588 2664
rect 4596 2656 4598 2664
rect 4586 2654 4598 2656
rect 4682 2764 4694 2766
rect 4682 2756 4684 2764
rect 4692 2756 4694 2764
rect 4682 2544 4694 2756
rect 4682 2536 4684 2544
rect 4692 2536 4694 2544
rect 4682 2534 4694 2536
rect 4522 2176 4524 2184
rect 4532 2176 4534 2184
rect 4522 2174 4534 2176
rect 4554 2524 4566 2526
rect 4554 2516 4556 2524
rect 4564 2516 4566 2524
rect 4416 2006 4420 2014
rect 4428 2006 4432 2014
rect 4440 2006 4444 2014
rect 4452 2006 4456 2014
rect 4464 2006 4468 2014
rect 4476 2006 4480 2014
rect 4416 1614 4480 2006
rect 4416 1606 4420 1614
rect 4428 1606 4432 1614
rect 4440 1606 4444 1614
rect 4452 1606 4456 1614
rect 4464 1606 4468 1614
rect 4476 1606 4480 1614
rect 4416 1214 4480 1606
rect 4416 1206 4420 1214
rect 4428 1206 4432 1214
rect 4440 1206 4444 1214
rect 4452 1206 4456 1214
rect 4464 1206 4468 1214
rect 4476 1206 4480 1214
rect 4330 736 4332 744
rect 4340 736 4342 744
rect 4330 734 4342 736
rect 4362 1124 4374 1126
rect 4362 1116 4364 1124
rect 4372 1116 4374 1124
rect 4362 524 4374 1116
rect 4362 516 4364 524
rect 4372 516 4374 524
rect 4362 514 4374 516
rect 4416 814 4480 1206
rect 4522 1884 4534 1886
rect 4522 1876 4524 1884
rect 4532 1876 4534 1884
rect 4522 1104 4534 1876
rect 4554 1644 4566 2516
rect 4586 2504 4598 2506
rect 4586 2496 4588 2504
rect 4596 2496 4598 2504
rect 4586 2324 4598 2496
rect 4714 2464 4726 2896
rect 5226 2604 5238 2606
rect 5226 2596 5228 2604
rect 5236 2596 5238 2604
rect 5226 2524 5238 2596
rect 5226 2516 5228 2524
rect 5236 2516 5238 2524
rect 5226 2514 5238 2516
rect 5546 2544 5558 2546
rect 5546 2536 5548 2544
rect 5556 2536 5558 2544
rect 4714 2456 4716 2464
rect 4724 2456 4726 2464
rect 4714 2454 4726 2456
rect 4842 2504 4854 2506
rect 4842 2496 4844 2504
rect 4852 2496 4854 2504
rect 4586 2316 4588 2324
rect 4596 2316 4598 2324
rect 4586 2314 4598 2316
rect 4746 2324 4758 2326
rect 4746 2316 4748 2324
rect 4756 2316 4758 2324
rect 4714 2304 4726 2306
rect 4714 2296 4716 2304
rect 4724 2296 4726 2304
rect 4586 2284 4598 2286
rect 4586 2276 4588 2284
rect 4596 2276 4598 2284
rect 4586 1724 4598 2276
rect 4650 2284 4662 2286
rect 4650 2276 4652 2284
rect 4660 2276 4662 2284
rect 4650 2124 4662 2276
rect 4650 2116 4652 2124
rect 4660 2116 4662 2124
rect 4650 2114 4662 2116
rect 4714 2124 4726 2296
rect 4714 2116 4716 2124
rect 4724 2116 4726 2124
rect 4714 2114 4726 2116
rect 4586 1716 4588 1724
rect 4596 1716 4598 1724
rect 4586 1714 4598 1716
rect 4682 2084 4694 2086
rect 4682 2076 4684 2084
rect 4692 2076 4694 2084
rect 4554 1636 4556 1644
rect 4564 1636 4566 1644
rect 4554 1634 4566 1636
rect 4586 1484 4598 1486
rect 4586 1476 4588 1484
rect 4596 1476 4598 1484
rect 4554 1324 4566 1326
rect 4554 1316 4556 1324
rect 4564 1316 4566 1324
rect 4554 1244 4566 1316
rect 4554 1236 4556 1244
rect 4564 1236 4566 1244
rect 4554 1234 4566 1236
rect 4522 1096 4524 1104
rect 4532 1096 4534 1104
rect 4522 1094 4534 1096
rect 4416 806 4420 814
rect 4428 806 4432 814
rect 4440 806 4444 814
rect 4452 806 4456 814
rect 4464 806 4468 814
rect 4476 806 4480 814
rect 4298 356 4300 364
rect 4308 356 4310 364
rect 4042 276 4044 284
rect 4052 276 4054 284
rect 4042 274 4054 276
rect 4074 304 4086 306
rect 4074 296 4076 304
rect 4084 296 4086 304
rect 3882 176 3884 184
rect 3892 176 3894 184
rect 3882 174 3894 176
rect 3754 96 3756 104
rect 3764 96 3766 104
rect 3754 94 3766 96
rect 3658 16 3660 24
rect 3668 16 3670 24
rect 3658 14 3670 16
rect 4074 24 4086 296
rect 4298 284 4310 356
rect 4298 276 4300 284
rect 4308 276 4310 284
rect 4298 274 4310 276
rect 4416 414 4480 806
rect 4522 1064 4534 1066
rect 4522 1056 4524 1064
rect 4532 1056 4534 1064
rect 4522 584 4534 1056
rect 4586 884 4598 1476
rect 4650 1484 4662 1486
rect 4650 1476 4652 1484
rect 4660 1476 4662 1484
rect 4650 1304 4662 1476
rect 4682 1384 4694 2076
rect 4746 1484 4758 2316
rect 4842 2284 4854 2496
rect 5482 2444 5494 2446
rect 5482 2436 5484 2444
rect 5492 2436 5494 2444
rect 5482 2364 5494 2436
rect 5482 2356 5484 2364
rect 5492 2356 5494 2364
rect 5482 2354 5494 2356
rect 4842 2276 4844 2284
rect 4852 2276 4854 2284
rect 4842 2274 4854 2276
rect 5066 2304 5078 2306
rect 5066 2296 5068 2304
rect 5076 2296 5078 2304
rect 4970 2184 4982 2186
rect 4970 2176 4972 2184
rect 4980 2176 4982 2184
rect 4970 1844 4982 2176
rect 4970 1836 4972 1844
rect 4980 1836 4982 1844
rect 4970 1834 4982 1836
rect 5002 2164 5014 2166
rect 5002 2156 5004 2164
rect 5012 2156 5014 2164
rect 4746 1476 4748 1484
rect 4756 1476 4758 1484
rect 4746 1474 4758 1476
rect 4810 1704 4822 1706
rect 4810 1696 4812 1704
rect 4820 1696 4822 1704
rect 4682 1376 4684 1384
rect 4692 1376 4694 1384
rect 4682 1374 4694 1376
rect 4650 1296 4652 1304
rect 4660 1296 4662 1304
rect 4650 1294 4662 1296
rect 4586 876 4588 884
rect 4596 876 4598 884
rect 4586 874 4598 876
rect 4618 1084 4630 1086
rect 4618 1076 4620 1084
rect 4628 1076 4630 1084
rect 4522 576 4524 584
rect 4532 576 4534 584
rect 4522 574 4534 576
rect 4416 406 4420 414
rect 4428 406 4432 414
rect 4440 406 4444 414
rect 4452 406 4456 414
rect 4464 406 4468 414
rect 4476 406 4480 414
rect 4074 16 4076 24
rect 4084 16 4086 24
rect 4074 14 4086 16
rect 4416 14 4480 406
rect 4618 284 4630 1076
rect 4778 924 4790 926
rect 4778 916 4780 924
rect 4788 916 4790 924
rect 4746 904 4758 906
rect 4746 896 4748 904
rect 4756 896 4758 904
rect 4618 276 4620 284
rect 4628 276 4630 284
rect 4618 184 4630 276
rect 4618 176 4620 184
rect 4628 176 4630 184
rect 4618 174 4630 176
rect 4650 544 4662 546
rect 4650 536 4652 544
rect 4660 536 4662 544
rect 4650 144 4662 536
rect 4746 524 4758 896
rect 4778 684 4790 916
rect 4778 676 4780 684
rect 4788 676 4790 684
rect 4778 674 4790 676
rect 4810 584 4822 1696
rect 4938 1644 4950 1646
rect 4938 1636 4940 1644
rect 4948 1636 4950 1644
rect 4938 1604 4950 1636
rect 4938 1596 4940 1604
rect 4948 1596 4950 1604
rect 4938 1594 4950 1596
rect 4874 1484 4886 1486
rect 4874 1476 4876 1484
rect 4884 1476 4886 1484
rect 4810 576 4812 584
rect 4820 576 4822 584
rect 4810 574 4822 576
rect 4842 804 4854 806
rect 4842 796 4844 804
rect 4852 796 4854 804
rect 4746 516 4748 524
rect 4756 516 4758 524
rect 4746 514 4758 516
rect 4650 136 4652 144
rect 4660 136 4662 144
rect 4650 134 4662 136
rect 4810 304 4822 306
rect 4810 296 4812 304
rect 4820 296 4822 304
rect 4810 44 4822 296
rect 4842 304 4854 796
rect 4874 784 4886 1476
rect 4938 1464 4950 1466
rect 4938 1456 4940 1464
rect 4948 1456 4950 1464
rect 4938 1364 4950 1456
rect 4938 1356 4940 1364
rect 4948 1356 4950 1364
rect 4938 1354 4950 1356
rect 4970 1424 4982 1426
rect 4970 1416 4972 1424
rect 4980 1416 4982 1424
rect 4874 776 4876 784
rect 4884 776 4886 784
rect 4874 774 4886 776
rect 4906 1124 4918 1126
rect 4906 1116 4908 1124
rect 4916 1116 4918 1124
rect 4842 296 4844 304
rect 4852 296 4854 304
rect 4842 294 4854 296
rect 4874 684 4886 686
rect 4874 676 4876 684
rect 4884 676 4886 684
rect 4842 204 4854 206
rect 4842 196 4844 204
rect 4852 196 4854 204
rect 4842 104 4854 196
rect 4842 96 4844 104
rect 4852 96 4854 104
rect 4842 94 4854 96
rect 4874 84 4886 676
rect 4906 524 4918 1116
rect 4906 516 4908 524
rect 4916 516 4918 524
rect 4906 514 4918 516
rect 4938 724 4950 726
rect 4938 716 4940 724
rect 4948 716 4950 724
rect 4938 244 4950 716
rect 4970 624 4982 1416
rect 4970 616 4972 624
rect 4980 616 4982 624
rect 4970 614 4982 616
rect 5002 544 5014 2156
rect 5066 1824 5078 2296
rect 5066 1816 5068 1824
rect 5076 1816 5078 1824
rect 5066 1814 5078 1816
rect 5098 2024 5110 2026
rect 5098 2016 5100 2024
rect 5108 2016 5110 2024
rect 5098 1764 5110 2016
rect 5098 1756 5100 1764
rect 5108 1756 5110 1764
rect 5098 1754 5110 1756
rect 5130 1824 5142 1826
rect 5130 1816 5132 1824
rect 5140 1816 5142 1824
rect 5098 1284 5110 1286
rect 5098 1276 5100 1284
rect 5108 1276 5110 1284
rect 5066 1104 5078 1106
rect 5066 1096 5068 1104
rect 5076 1096 5078 1104
rect 5002 536 5004 544
rect 5012 536 5014 544
rect 5002 534 5014 536
rect 5034 664 5046 666
rect 5034 656 5036 664
rect 5044 656 5046 664
rect 4938 236 4940 244
rect 4948 236 4950 244
rect 4938 234 4950 236
rect 5034 164 5046 656
rect 5034 156 5036 164
rect 5044 156 5046 164
rect 5034 154 5046 156
rect 5066 104 5078 1096
rect 5098 284 5110 1276
rect 5130 1124 5142 1816
rect 5546 1764 5558 2536
rect 5578 2524 5590 2916
rect 5578 2516 5580 2524
rect 5588 2516 5590 2524
rect 5578 2514 5590 2516
rect 5642 2524 5654 4136
rect 5674 4104 5686 4106
rect 5674 4096 5676 4104
rect 5684 4096 5686 4104
rect 5674 3964 5686 4096
rect 5674 3956 5676 3964
rect 5684 3956 5686 3964
rect 5674 3954 5686 3956
rect 5738 3644 5750 4196
rect 5770 4144 5782 4296
rect 5770 4136 5772 4144
rect 5780 4136 5782 4144
rect 5770 4134 5782 4136
rect 5802 4304 5814 4676
rect 5802 4296 5804 4304
rect 5812 4296 5814 4304
rect 5802 4104 5814 4296
rect 5866 4304 5878 4696
rect 5866 4296 5868 4304
rect 5876 4296 5878 4304
rect 5802 4096 5804 4104
rect 5812 4096 5814 4104
rect 5802 4094 5814 4096
rect 5834 4164 5846 4166
rect 5834 4156 5836 4164
rect 5844 4156 5846 4164
rect 5834 4084 5846 4156
rect 5866 4124 5878 4296
rect 5866 4116 5868 4124
rect 5876 4116 5878 4124
rect 5866 4114 5878 4116
rect 5920 4614 5984 5006
rect 6186 5104 6198 5106
rect 6186 5096 6188 5104
rect 6196 5096 6198 5104
rect 5920 4606 5924 4614
rect 5932 4606 5936 4614
rect 5944 4606 5948 4614
rect 5956 4606 5960 4614
rect 5968 4606 5972 4614
rect 5980 4606 5984 4614
rect 5920 4214 5984 4606
rect 6026 4904 6038 4906
rect 6026 4896 6028 4904
rect 6036 4896 6038 4904
rect 6026 4564 6038 4896
rect 6186 4844 6198 5096
rect 6858 5104 6870 5106
rect 6858 5096 6860 5104
rect 6868 5096 6870 5104
rect 6186 4836 6188 4844
rect 6196 4836 6198 4844
rect 6186 4834 6198 4836
rect 6378 5024 6390 5026
rect 6378 5016 6380 5024
rect 6388 5016 6390 5024
rect 6058 4824 6070 4826
rect 6058 4816 6060 4824
rect 6068 4816 6070 4824
rect 6058 4704 6070 4816
rect 6058 4696 6060 4704
rect 6068 4696 6070 4704
rect 6058 4694 6070 4696
rect 6026 4556 6028 4564
rect 6036 4556 6038 4564
rect 6026 4554 6038 4556
rect 6122 4564 6134 4566
rect 6122 4556 6124 4564
rect 6132 4556 6134 4564
rect 6122 4384 6134 4556
rect 6314 4544 6326 4546
rect 6314 4536 6316 4544
rect 6324 4536 6326 4544
rect 6218 4524 6230 4526
rect 6218 4516 6220 4524
rect 6228 4516 6230 4524
rect 6186 4484 6198 4486
rect 6186 4476 6188 4484
rect 6196 4476 6198 4484
rect 6186 4424 6198 4476
rect 6186 4416 6188 4424
rect 6196 4416 6198 4424
rect 6122 4376 6124 4384
rect 6132 4376 6134 4384
rect 6122 4374 6134 4376
rect 6154 4384 6166 4386
rect 6154 4376 6156 4384
rect 6164 4376 6166 4384
rect 5920 4206 5924 4214
rect 5932 4206 5936 4214
rect 5944 4206 5948 4214
rect 5956 4206 5960 4214
rect 5968 4206 5972 4214
rect 5980 4206 5984 4214
rect 5834 4076 5836 4084
rect 5844 4076 5846 4084
rect 5834 4074 5846 4076
rect 5738 3636 5740 3644
rect 5748 3636 5750 3644
rect 5738 3634 5750 3636
rect 5770 3924 5782 3926
rect 5770 3916 5772 3924
rect 5780 3916 5782 3924
rect 5770 3884 5782 3916
rect 5770 3876 5772 3884
rect 5780 3876 5782 3884
rect 5770 3284 5782 3876
rect 5770 3276 5772 3284
rect 5780 3276 5782 3284
rect 5770 3204 5782 3276
rect 5770 3196 5772 3204
rect 5780 3196 5782 3204
rect 5770 3194 5782 3196
rect 5920 3814 5984 4206
rect 6122 4344 6134 4346
rect 6122 4336 6124 4344
rect 6132 4336 6134 4344
rect 5920 3806 5924 3814
rect 5932 3806 5936 3814
rect 5944 3806 5948 3814
rect 5956 3806 5960 3814
rect 5968 3806 5972 3814
rect 5980 3806 5984 3814
rect 5920 3414 5984 3806
rect 6058 3844 6070 3846
rect 6058 3836 6060 3844
rect 6068 3836 6070 3844
rect 6026 3564 6038 3566
rect 6026 3556 6028 3564
rect 6036 3556 6038 3564
rect 6026 3484 6038 3556
rect 6058 3504 6070 3836
rect 6058 3496 6060 3504
rect 6068 3496 6070 3504
rect 6058 3494 6070 3496
rect 6090 3664 6102 3666
rect 6090 3656 6092 3664
rect 6100 3656 6102 3664
rect 6026 3476 6028 3484
rect 6036 3476 6038 3484
rect 6026 3474 6038 3476
rect 5920 3406 5924 3414
rect 5932 3406 5936 3414
rect 5944 3406 5948 3414
rect 5956 3406 5960 3414
rect 5968 3406 5972 3414
rect 5980 3406 5984 3414
rect 5920 3014 5984 3406
rect 5920 3006 5924 3014
rect 5932 3006 5936 3014
rect 5944 3006 5948 3014
rect 5956 3006 5960 3014
rect 5968 3006 5972 3014
rect 5980 3006 5984 3014
rect 5834 2904 5846 2906
rect 5834 2896 5836 2904
rect 5844 2896 5846 2904
rect 5642 2516 5644 2524
rect 5652 2516 5654 2524
rect 5642 2514 5654 2516
rect 5738 2684 5750 2686
rect 5738 2676 5740 2684
rect 5748 2676 5750 2684
rect 5610 2504 5622 2506
rect 5610 2496 5612 2504
rect 5620 2496 5622 2504
rect 5610 2304 5622 2496
rect 5610 2296 5612 2304
rect 5620 2296 5622 2304
rect 5610 2294 5622 2296
rect 5642 2484 5654 2486
rect 5642 2476 5644 2484
rect 5652 2476 5654 2484
rect 5642 2284 5654 2476
rect 5738 2484 5750 2676
rect 5802 2664 5814 2666
rect 5802 2656 5804 2664
rect 5812 2656 5814 2664
rect 5802 2564 5814 2656
rect 5834 2624 5846 2896
rect 5834 2616 5836 2624
rect 5844 2616 5846 2624
rect 5834 2614 5846 2616
rect 5920 2614 5984 3006
rect 6026 3424 6038 3426
rect 6026 3416 6028 3424
rect 6036 3416 6038 3424
rect 6026 2684 6038 3416
rect 6090 3404 6102 3656
rect 6090 3396 6092 3404
rect 6100 3396 6102 3404
rect 6090 3394 6102 3396
rect 6122 3384 6134 4336
rect 6122 3376 6124 3384
rect 6132 3376 6134 3384
rect 6122 3374 6134 3376
rect 6154 3304 6166 4376
rect 6186 3524 6198 4416
rect 6218 4164 6230 4516
rect 6314 4504 6326 4536
rect 6314 4496 6316 4504
rect 6324 4496 6326 4504
rect 6314 4494 6326 4496
rect 6314 4404 6326 4406
rect 6314 4396 6316 4404
rect 6324 4396 6326 4404
rect 6218 4156 6220 4164
rect 6228 4156 6230 4164
rect 6218 4154 6230 4156
rect 6250 4304 6262 4306
rect 6250 4296 6252 4304
rect 6260 4296 6262 4304
rect 6250 4124 6262 4296
rect 6250 4116 6252 4124
rect 6260 4116 6262 4124
rect 6250 4114 6262 4116
rect 6282 4184 6294 4186
rect 6282 4176 6284 4184
rect 6292 4176 6294 4184
rect 6250 3864 6262 3866
rect 6250 3856 6252 3864
rect 6260 3856 6262 3864
rect 6186 3516 6188 3524
rect 6196 3516 6198 3524
rect 6186 3514 6198 3516
rect 6218 3644 6230 3646
rect 6218 3636 6220 3644
rect 6228 3636 6230 3644
rect 6154 3296 6156 3304
rect 6164 3296 6166 3304
rect 6154 3294 6166 3296
rect 6186 3404 6198 3406
rect 6186 3396 6188 3404
rect 6196 3396 6198 3404
rect 6186 3084 6198 3396
rect 6186 3076 6188 3084
rect 6196 3076 6198 3084
rect 6186 3074 6198 3076
rect 6218 2924 6230 3636
rect 6250 2944 6262 3856
rect 6282 3864 6294 4176
rect 6314 4184 6326 4396
rect 6314 4176 6316 4184
rect 6324 4176 6326 4184
rect 6314 4174 6326 4176
rect 6282 3856 6284 3864
rect 6292 3856 6294 3864
rect 6282 3854 6294 3856
rect 6346 3104 6358 3106
rect 6346 3096 6348 3104
rect 6356 3096 6358 3104
rect 6282 3084 6294 3086
rect 6282 3076 6284 3084
rect 6292 3076 6294 3084
rect 6282 2964 6294 3076
rect 6282 2956 6284 2964
rect 6292 2956 6294 2964
rect 6282 2954 6294 2956
rect 6250 2936 6252 2944
rect 6260 2936 6262 2944
rect 6250 2934 6262 2936
rect 6218 2916 6220 2924
rect 6228 2916 6230 2924
rect 6218 2914 6230 2916
rect 6026 2676 6028 2684
rect 6036 2676 6038 2684
rect 6026 2674 6038 2676
rect 6282 2684 6294 2686
rect 6282 2676 6284 2684
rect 6292 2676 6294 2684
rect 5802 2556 5804 2564
rect 5812 2556 5814 2564
rect 5802 2554 5814 2556
rect 5920 2606 5924 2614
rect 5932 2606 5936 2614
rect 5944 2606 5948 2614
rect 5956 2606 5960 2614
rect 5968 2606 5972 2614
rect 5980 2606 5984 2614
rect 5738 2476 5740 2484
rect 5748 2476 5750 2484
rect 5738 2474 5750 2476
rect 5642 2276 5644 2284
rect 5652 2276 5654 2284
rect 5578 1984 5590 1986
rect 5578 1976 5580 1984
rect 5588 1976 5590 1984
rect 5578 1784 5590 1976
rect 5578 1776 5580 1784
rect 5588 1776 5590 1784
rect 5578 1774 5590 1776
rect 5546 1756 5548 1764
rect 5556 1756 5558 1764
rect 5546 1754 5558 1756
rect 5194 1664 5206 1666
rect 5194 1656 5196 1664
rect 5204 1656 5206 1664
rect 5194 1264 5206 1656
rect 5322 1604 5334 1606
rect 5322 1596 5324 1604
rect 5332 1596 5334 1604
rect 5258 1544 5270 1546
rect 5258 1536 5260 1544
rect 5268 1536 5270 1544
rect 5258 1464 5270 1536
rect 5258 1456 5260 1464
rect 5268 1456 5270 1464
rect 5258 1454 5270 1456
rect 5290 1484 5302 1486
rect 5290 1476 5292 1484
rect 5300 1476 5302 1484
rect 5290 1304 5302 1476
rect 5290 1296 5292 1304
rect 5300 1296 5302 1304
rect 5290 1294 5302 1296
rect 5194 1256 5196 1264
rect 5204 1256 5206 1264
rect 5194 1144 5206 1256
rect 5194 1136 5196 1144
rect 5204 1136 5206 1144
rect 5194 1134 5206 1136
rect 5130 1116 5132 1124
rect 5140 1116 5142 1124
rect 5130 1114 5142 1116
rect 5322 1104 5334 1596
rect 5610 1524 5622 1526
rect 5610 1516 5612 1524
rect 5620 1516 5622 1524
rect 5546 1504 5558 1506
rect 5546 1496 5548 1504
rect 5556 1496 5558 1504
rect 5322 1096 5324 1104
rect 5332 1096 5334 1104
rect 5322 1094 5334 1096
rect 5450 1404 5462 1406
rect 5450 1396 5452 1404
rect 5460 1396 5462 1404
rect 5450 1144 5462 1396
rect 5546 1384 5558 1496
rect 5610 1464 5622 1516
rect 5610 1456 5612 1464
rect 5620 1456 5622 1464
rect 5610 1454 5622 1456
rect 5642 1424 5654 2276
rect 5706 2364 5718 2366
rect 5706 2356 5708 2364
rect 5716 2356 5718 2364
rect 5706 2224 5718 2356
rect 5706 2216 5708 2224
rect 5716 2216 5718 2224
rect 5706 2214 5718 2216
rect 5802 2324 5814 2326
rect 5802 2316 5804 2324
rect 5812 2316 5814 2324
rect 5770 1884 5782 1886
rect 5770 1876 5772 1884
rect 5780 1876 5782 1884
rect 5770 1624 5782 1876
rect 5770 1616 5772 1624
rect 5780 1616 5782 1624
rect 5770 1614 5782 1616
rect 5642 1416 5644 1424
rect 5652 1416 5654 1424
rect 5642 1414 5654 1416
rect 5546 1376 5548 1384
rect 5556 1376 5558 1384
rect 5546 1374 5558 1376
rect 5450 1136 5452 1144
rect 5460 1136 5462 1144
rect 5450 944 5462 1136
rect 5450 936 5452 944
rect 5460 936 5462 944
rect 5450 934 5462 936
rect 5610 1084 5622 1086
rect 5610 1076 5612 1084
rect 5620 1076 5622 1084
rect 5098 276 5100 284
rect 5108 276 5110 284
rect 5098 274 5110 276
rect 5194 604 5206 606
rect 5194 596 5196 604
rect 5204 596 5206 604
rect 5066 96 5068 104
rect 5076 96 5078 104
rect 5066 94 5078 96
rect 4874 76 4876 84
rect 4884 76 4886 84
rect 4874 74 4886 76
rect 4810 36 4812 44
rect 4820 36 4822 44
rect 4810 34 4822 36
rect 5194 24 5206 596
rect 5610 604 5622 1076
rect 5770 924 5782 926
rect 5770 916 5772 924
rect 5780 916 5782 924
rect 5770 624 5782 916
rect 5802 904 5814 2316
rect 5802 896 5804 904
rect 5812 896 5814 904
rect 5802 724 5814 896
rect 5802 716 5804 724
rect 5812 716 5814 724
rect 5802 714 5814 716
rect 5920 2214 5984 2606
rect 5920 2206 5924 2214
rect 5932 2206 5936 2214
rect 5944 2206 5948 2214
rect 5956 2206 5960 2214
rect 5968 2206 5972 2214
rect 5980 2206 5984 2214
rect 5920 1814 5984 2206
rect 6026 2524 6038 2526
rect 6026 2516 6028 2524
rect 6036 2516 6038 2524
rect 6026 1844 6038 2516
rect 6282 2324 6294 2676
rect 6282 2316 6284 2324
rect 6292 2316 6294 2324
rect 6282 2314 6294 2316
rect 6154 2304 6166 2306
rect 6154 2296 6156 2304
rect 6164 2296 6166 2304
rect 6154 2084 6166 2296
rect 6218 2224 6230 2226
rect 6218 2216 6220 2224
rect 6228 2216 6230 2224
rect 6218 2164 6230 2216
rect 6218 2156 6220 2164
rect 6228 2156 6230 2164
rect 6218 2154 6230 2156
rect 6314 2184 6326 2186
rect 6314 2176 6316 2184
rect 6324 2176 6326 2184
rect 6154 2076 6156 2084
rect 6164 2076 6166 2084
rect 6154 2074 6166 2076
rect 6154 2044 6166 2046
rect 6154 2036 6156 2044
rect 6164 2036 6166 2044
rect 6026 1836 6028 1844
rect 6036 1836 6038 1844
rect 6026 1834 6038 1836
rect 6058 1904 6070 1906
rect 6058 1896 6060 1904
rect 6068 1896 6070 1904
rect 5920 1806 5924 1814
rect 5932 1806 5936 1814
rect 5944 1806 5948 1814
rect 5956 1806 5960 1814
rect 5968 1806 5972 1814
rect 5980 1806 5984 1814
rect 5920 1414 5984 1806
rect 5920 1406 5924 1414
rect 5932 1406 5936 1414
rect 5944 1406 5948 1414
rect 5956 1406 5960 1414
rect 5968 1406 5972 1414
rect 5980 1406 5984 1414
rect 5920 1014 5984 1406
rect 6026 1564 6038 1566
rect 6026 1556 6028 1564
rect 6036 1556 6038 1564
rect 6026 1264 6038 1556
rect 6026 1256 6028 1264
rect 6036 1256 6038 1264
rect 6026 1254 6038 1256
rect 5920 1006 5924 1014
rect 5932 1006 5936 1014
rect 5944 1006 5948 1014
rect 5956 1006 5960 1014
rect 5968 1006 5972 1014
rect 5980 1006 5984 1014
rect 5770 616 5772 624
rect 5780 616 5782 624
rect 5770 614 5782 616
rect 5920 614 5984 1006
rect 6026 1024 6038 1026
rect 6026 1016 6028 1024
rect 6036 1016 6038 1024
rect 6026 704 6038 1016
rect 6026 696 6028 704
rect 6036 696 6038 704
rect 6026 694 6038 696
rect 5610 596 5612 604
rect 5620 596 5622 604
rect 5610 594 5622 596
rect 5920 606 5924 614
rect 5932 606 5936 614
rect 5944 606 5948 614
rect 5956 606 5960 614
rect 5968 606 5972 614
rect 5980 606 5984 614
rect 5802 524 5814 526
rect 5802 516 5804 524
rect 5812 516 5814 524
rect 5802 464 5814 516
rect 5802 456 5804 464
rect 5812 456 5814 464
rect 5802 454 5814 456
rect 5194 16 5196 24
rect 5204 16 5206 24
rect 5194 14 5206 16
rect 5920 214 5984 606
rect 6058 484 6070 1896
rect 6154 1884 6166 2036
rect 6154 1876 6156 1884
rect 6164 1876 6166 1884
rect 6154 1874 6166 1876
rect 6282 2024 6294 2026
rect 6282 2016 6284 2024
rect 6292 2016 6294 2024
rect 6090 1864 6102 1866
rect 6090 1856 6092 1864
rect 6100 1856 6102 1864
rect 6090 1284 6102 1856
rect 6282 1784 6294 2016
rect 6314 1864 6326 2176
rect 6346 2144 6358 3096
rect 6346 2136 6348 2144
rect 6356 2136 6358 2144
rect 6346 2134 6358 2136
rect 6314 1856 6316 1864
rect 6324 1856 6326 1864
rect 6314 1854 6326 1856
rect 6282 1776 6284 1784
rect 6292 1776 6294 1784
rect 6282 1774 6294 1776
rect 6314 1784 6326 1786
rect 6314 1776 6316 1784
rect 6324 1776 6326 1784
rect 6186 1744 6198 1746
rect 6186 1736 6188 1744
rect 6196 1736 6198 1744
rect 6090 1276 6092 1284
rect 6100 1276 6102 1284
rect 6090 1274 6102 1276
rect 6122 1724 6134 1726
rect 6122 1716 6124 1724
rect 6132 1716 6134 1724
rect 6122 584 6134 1716
rect 6186 1244 6198 1736
rect 6314 1704 6326 1776
rect 6314 1696 6316 1704
rect 6324 1696 6326 1704
rect 6314 1694 6326 1696
rect 6218 1584 6230 1586
rect 6218 1576 6220 1584
rect 6228 1576 6230 1584
rect 6218 1344 6230 1576
rect 6218 1336 6220 1344
rect 6228 1336 6230 1344
rect 6218 1334 6230 1336
rect 6282 1464 6294 1466
rect 6282 1456 6284 1464
rect 6292 1456 6294 1464
rect 6186 1236 6188 1244
rect 6196 1236 6198 1244
rect 6186 1104 6198 1236
rect 6186 1096 6188 1104
rect 6196 1096 6198 1104
rect 6186 1094 6198 1096
rect 6250 1304 6262 1306
rect 6250 1296 6252 1304
rect 6260 1296 6262 1304
rect 6122 576 6124 584
rect 6132 576 6134 584
rect 6122 574 6134 576
rect 6186 1044 6198 1046
rect 6186 1036 6188 1044
rect 6196 1036 6198 1044
rect 6058 476 6060 484
rect 6068 476 6070 484
rect 6058 474 6070 476
rect 6186 324 6198 1036
rect 6250 904 6262 1296
rect 6282 1144 6294 1456
rect 6282 1136 6284 1144
rect 6292 1136 6294 1144
rect 6282 1134 6294 1136
rect 6250 896 6252 904
rect 6260 896 6262 904
rect 6250 894 6262 896
rect 6282 744 6294 746
rect 6282 736 6284 744
rect 6292 736 6294 744
rect 6282 704 6294 736
rect 6282 696 6284 704
rect 6292 696 6294 704
rect 6282 694 6294 696
rect 6186 316 6188 324
rect 6196 316 6198 324
rect 6186 314 6198 316
rect 5920 206 5924 214
rect 5932 206 5936 214
rect 5944 206 5948 214
rect 5956 206 5960 214
rect 5968 206 5972 214
rect 5980 206 5984 214
rect 4416 6 4420 14
rect 4428 6 4432 14
rect 4440 6 4444 14
rect 4452 6 4456 14
rect 4464 6 4468 14
rect 4476 6 4480 14
rect 4416 -10 4480 6
rect 5920 -10 5984 206
rect 6378 164 6390 5016
rect 6570 4704 6582 4706
rect 6570 4696 6572 4704
rect 6580 4696 6582 4704
rect 6570 4544 6582 4696
rect 6570 4536 6572 4544
rect 6580 4536 6582 4544
rect 6570 4284 6582 4536
rect 6570 4276 6572 4284
rect 6580 4276 6582 4284
rect 6570 4274 6582 4276
rect 6442 4064 6454 4066
rect 6442 4056 6444 4064
rect 6452 4056 6454 4064
rect 6442 3844 6454 4056
rect 6570 4024 6582 4026
rect 6570 4016 6572 4024
rect 6580 4016 6582 4024
rect 6442 3836 6444 3844
rect 6452 3836 6454 3844
rect 6442 3834 6454 3836
rect 6474 3884 6486 3886
rect 6474 3876 6476 3884
rect 6484 3876 6486 3884
rect 6474 3784 6486 3876
rect 6474 3776 6476 3784
rect 6484 3776 6486 3784
rect 6442 3704 6454 3706
rect 6442 3696 6444 3704
rect 6452 3696 6454 3704
rect 6442 2524 6454 3696
rect 6474 3504 6486 3776
rect 6570 3584 6582 4016
rect 6698 4004 6710 4006
rect 6698 3996 6700 4004
rect 6708 3996 6710 4004
rect 6570 3576 6572 3584
rect 6580 3576 6582 3584
rect 6570 3574 6582 3576
rect 6666 3984 6678 3986
rect 6666 3976 6668 3984
rect 6676 3976 6678 3984
rect 6666 3564 6678 3976
rect 6698 3644 6710 3996
rect 6698 3636 6700 3644
rect 6708 3636 6710 3644
rect 6698 3634 6710 3636
rect 6730 3684 6742 3686
rect 6730 3676 6732 3684
rect 6740 3676 6742 3684
rect 6666 3556 6668 3564
rect 6676 3556 6678 3564
rect 6666 3554 6678 3556
rect 6474 3496 6476 3504
rect 6484 3496 6486 3504
rect 6474 3494 6486 3496
rect 6634 3324 6646 3326
rect 6634 3316 6636 3324
rect 6644 3316 6646 3324
rect 6442 2516 6444 2524
rect 6452 2516 6454 2524
rect 6442 2514 6454 2516
rect 6474 2964 6486 2966
rect 6474 2956 6476 2964
rect 6484 2956 6486 2964
rect 6410 1964 6422 1966
rect 6410 1956 6412 1964
rect 6420 1956 6422 1964
rect 6410 1824 6422 1956
rect 6410 1816 6412 1824
rect 6420 1816 6422 1824
rect 6410 1814 6422 1816
rect 6442 1824 6454 1826
rect 6442 1816 6444 1824
rect 6452 1816 6454 1824
rect 6442 1744 6454 1816
rect 6442 1736 6444 1744
rect 6452 1736 6454 1744
rect 6442 1734 6454 1736
rect 6474 1584 6486 2956
rect 6570 2304 6582 2306
rect 6570 2296 6572 2304
rect 6580 2296 6582 2304
rect 6570 1884 6582 2296
rect 6570 1876 6572 1884
rect 6580 1876 6582 1884
rect 6570 1724 6582 1876
rect 6570 1716 6572 1724
rect 6580 1716 6582 1724
rect 6570 1714 6582 1716
rect 6474 1576 6476 1584
rect 6484 1576 6486 1584
rect 6474 1574 6486 1576
rect 6602 1704 6614 1706
rect 6602 1696 6604 1704
rect 6612 1696 6614 1704
rect 6474 1544 6486 1546
rect 6474 1536 6476 1544
rect 6484 1536 6486 1544
rect 6442 1464 6454 1466
rect 6442 1456 6444 1464
rect 6452 1456 6454 1464
rect 6442 864 6454 1456
rect 6474 1424 6486 1536
rect 6474 1416 6476 1424
rect 6484 1416 6486 1424
rect 6474 1384 6486 1416
rect 6474 1376 6476 1384
rect 6484 1376 6486 1384
rect 6474 1374 6486 1376
rect 6602 1364 6614 1696
rect 6602 1356 6604 1364
rect 6612 1356 6614 1364
rect 6602 1354 6614 1356
rect 6602 1304 6614 1306
rect 6602 1296 6604 1304
rect 6612 1296 6614 1304
rect 6442 856 6444 864
rect 6452 856 6454 864
rect 6442 854 6454 856
rect 6474 1124 6486 1126
rect 6474 1116 6476 1124
rect 6484 1116 6486 1124
rect 6474 504 6486 1116
rect 6602 644 6614 1296
rect 6602 636 6604 644
rect 6612 636 6614 644
rect 6602 634 6614 636
rect 6474 496 6476 504
rect 6484 496 6486 504
rect 6474 494 6486 496
rect 6378 156 6380 164
rect 6388 156 6390 164
rect 6378 154 6390 156
rect 6634 104 6646 3316
rect 6730 2584 6742 3676
rect 6762 3644 6774 3646
rect 6762 3636 6764 3644
rect 6772 3636 6774 3644
rect 6762 3604 6774 3636
rect 6762 3596 6764 3604
rect 6772 3596 6774 3604
rect 6762 2744 6774 3596
rect 6826 3024 6838 3026
rect 6826 3016 6828 3024
rect 6836 3016 6838 3024
rect 6826 2964 6838 3016
rect 6826 2956 6828 2964
rect 6836 2956 6838 2964
rect 6826 2954 6838 2956
rect 6762 2736 6764 2744
rect 6772 2736 6774 2744
rect 6762 2734 6774 2736
rect 6794 2884 6806 2886
rect 6794 2876 6796 2884
rect 6804 2876 6806 2884
rect 6730 2576 6732 2584
rect 6740 2576 6742 2584
rect 6730 2574 6742 2576
rect 6698 2444 6710 2446
rect 6698 2436 6700 2444
rect 6708 2436 6710 2444
rect 6666 2204 6678 2206
rect 6666 2196 6668 2204
rect 6676 2196 6678 2204
rect 6666 1824 6678 2196
rect 6666 1816 6668 1824
rect 6676 1816 6678 1824
rect 6666 1814 6678 1816
rect 6698 1604 6710 2436
rect 6762 2344 6774 2346
rect 6762 2336 6764 2344
rect 6772 2336 6774 2344
rect 6698 1596 6700 1604
rect 6708 1596 6710 1604
rect 6698 1594 6710 1596
rect 6730 1824 6742 1826
rect 6730 1816 6732 1824
rect 6740 1816 6742 1824
rect 6666 844 6678 846
rect 6666 836 6668 844
rect 6676 836 6678 844
rect 6666 184 6678 836
rect 6698 784 6710 786
rect 6698 776 6700 784
rect 6708 776 6710 784
rect 6698 704 6710 776
rect 6698 696 6700 704
rect 6708 696 6710 704
rect 6698 694 6710 696
rect 6666 176 6668 184
rect 6676 176 6678 184
rect 6666 174 6678 176
rect 6730 184 6742 1816
rect 6762 1764 6774 2336
rect 6762 1756 6764 1764
rect 6772 1756 6774 1764
rect 6762 1754 6774 1756
rect 6794 1604 6806 2876
rect 6858 2524 6870 5096
rect 7370 5084 7382 5086
rect 7370 5076 7372 5084
rect 7380 5076 7382 5084
rect 7114 5044 7126 5046
rect 7114 5036 7116 5044
rect 7124 5036 7126 5044
rect 6954 4944 6966 4946
rect 6954 4936 6956 4944
rect 6964 4936 6966 4944
rect 6922 4524 6934 4526
rect 6922 4516 6924 4524
rect 6932 4516 6934 4524
rect 6890 3904 6902 3906
rect 6890 3896 6892 3904
rect 6900 3896 6902 3904
rect 6890 3504 6902 3896
rect 6890 3496 6892 3504
rect 6900 3496 6902 3504
rect 6890 3494 6902 3496
rect 6922 3124 6934 4516
rect 6954 3824 6966 4936
rect 7114 4904 7126 5036
rect 7114 4896 7116 4904
rect 7124 4896 7126 4904
rect 7082 4604 7094 4606
rect 7082 4596 7084 4604
rect 7092 4596 7094 4604
rect 6954 3816 6956 3824
rect 6964 3816 6966 3824
rect 6954 3814 6966 3816
rect 7018 3884 7030 3886
rect 7018 3876 7020 3884
rect 7028 3876 7030 3884
rect 6922 3116 6924 3124
rect 6932 3116 6934 3124
rect 6922 3114 6934 3116
rect 6954 3724 6966 3726
rect 6954 3716 6956 3724
rect 6964 3716 6966 3724
rect 6954 3084 6966 3716
rect 6986 3704 6998 3706
rect 6986 3696 6988 3704
rect 6996 3696 6998 3704
rect 6986 3344 6998 3696
rect 6986 3336 6988 3344
rect 6996 3336 6998 3344
rect 6986 3144 6998 3336
rect 6986 3136 6988 3144
rect 6996 3136 6998 3144
rect 6986 3134 6998 3136
rect 6954 3076 6956 3084
rect 6964 3076 6966 3084
rect 6954 3074 6966 3076
rect 6858 2516 6860 2524
rect 6868 2516 6870 2524
rect 6858 2514 6870 2516
rect 6922 3064 6934 3066
rect 6922 3056 6924 3064
rect 6932 3056 6934 3064
rect 6922 2184 6934 3056
rect 6922 2176 6924 2184
rect 6932 2176 6934 2184
rect 6922 2174 6934 2176
rect 6954 2484 6966 2486
rect 6954 2476 6956 2484
rect 6964 2476 6966 2484
rect 6954 2144 6966 2476
rect 6954 2136 6956 2144
rect 6964 2136 6966 2144
rect 6954 2134 6966 2136
rect 6986 2204 6998 2206
rect 6986 2196 6988 2204
rect 6996 2196 6998 2204
rect 6858 2124 6870 2126
rect 6858 2116 6860 2124
rect 6868 2116 6870 2124
rect 6794 1596 6796 1604
rect 6804 1596 6806 1604
rect 6794 1594 6806 1596
rect 6826 2044 6838 2046
rect 6826 2036 6828 2044
rect 6836 2036 6838 2044
rect 6826 1724 6838 2036
rect 6826 1716 6828 1724
rect 6836 1716 6838 1724
rect 6826 1344 6838 1716
rect 6858 1524 6870 2116
rect 6922 1924 6934 1926
rect 6922 1916 6924 1924
rect 6932 1916 6934 1924
rect 6858 1516 6860 1524
rect 6868 1516 6870 1524
rect 6858 1514 6870 1516
rect 6890 1904 6902 1906
rect 6890 1896 6892 1904
rect 6900 1896 6902 1904
rect 6826 1336 6828 1344
rect 6836 1336 6838 1344
rect 6826 1334 6838 1336
rect 6794 1324 6806 1326
rect 6794 1316 6796 1324
rect 6804 1316 6806 1324
rect 6794 304 6806 1316
rect 6890 1324 6902 1896
rect 6922 1444 6934 1916
rect 6986 1904 6998 2196
rect 6986 1896 6988 1904
rect 6996 1896 6998 1904
rect 6986 1894 6998 1896
rect 6954 1844 6966 1846
rect 6954 1836 6956 1844
rect 6964 1836 6966 1844
rect 6954 1724 6966 1836
rect 6954 1716 6956 1724
rect 6964 1716 6966 1724
rect 6954 1714 6966 1716
rect 6922 1436 6924 1444
rect 6932 1436 6934 1444
rect 6922 1434 6934 1436
rect 6954 1544 6966 1546
rect 6954 1536 6956 1544
rect 6964 1536 6966 1544
rect 6890 1316 6892 1324
rect 6900 1316 6902 1324
rect 6890 1314 6902 1316
rect 6922 1344 6934 1346
rect 6922 1336 6924 1344
rect 6932 1336 6934 1344
rect 6794 296 6796 304
rect 6804 296 6806 304
rect 6794 294 6806 296
rect 6730 176 6732 184
rect 6740 176 6742 184
rect 6730 174 6742 176
rect 6922 184 6934 1336
rect 6954 1124 6966 1536
rect 6954 1116 6956 1124
rect 6964 1116 6966 1124
rect 6954 1114 6966 1116
rect 6922 176 6924 184
rect 6932 176 6934 184
rect 6922 174 6934 176
rect 7018 144 7030 3876
rect 7082 3824 7094 4596
rect 7114 4524 7126 4896
rect 7306 5044 7318 5046
rect 7306 5036 7308 5044
rect 7316 5036 7318 5044
rect 7114 4516 7116 4524
rect 7124 4516 7126 4524
rect 7114 4514 7126 4516
rect 7146 4744 7158 4746
rect 7146 4736 7148 4744
rect 7156 4736 7158 4744
rect 7146 4324 7158 4736
rect 7274 4604 7286 4606
rect 7274 4596 7276 4604
rect 7284 4596 7286 4604
rect 7146 4316 7148 4324
rect 7156 4316 7158 4324
rect 7146 4314 7158 4316
rect 7210 4504 7222 4506
rect 7210 4496 7212 4504
rect 7220 4496 7222 4504
rect 7082 3816 7084 3824
rect 7092 3816 7094 3824
rect 7082 3814 7094 3816
rect 7146 4064 7158 4066
rect 7146 4056 7148 4064
rect 7156 4056 7158 4064
rect 7082 3744 7094 3746
rect 7082 3736 7084 3744
rect 7092 3736 7094 3744
rect 7050 3584 7062 3586
rect 7050 3576 7052 3584
rect 7060 3576 7062 3584
rect 7050 3104 7062 3576
rect 7082 3264 7094 3736
rect 7146 3364 7158 4056
rect 7146 3356 7148 3364
rect 7156 3356 7158 3364
rect 7146 3354 7158 3356
rect 7082 3256 7084 3264
rect 7092 3256 7094 3264
rect 7082 3254 7094 3256
rect 7210 3264 7222 4496
rect 7242 4124 7254 4126
rect 7242 4116 7244 4124
rect 7252 4116 7254 4124
rect 7242 3844 7254 4116
rect 7242 3836 7244 3844
rect 7252 3836 7254 3844
rect 7242 3834 7254 3836
rect 7210 3256 7212 3264
rect 7220 3256 7222 3264
rect 7210 3254 7222 3256
rect 7242 3764 7254 3766
rect 7242 3756 7244 3764
rect 7252 3756 7254 3764
rect 7050 3096 7052 3104
rect 7060 3096 7062 3104
rect 7050 3094 7062 3096
rect 7050 2984 7062 2986
rect 7050 2976 7052 2984
rect 7060 2976 7062 2984
rect 7050 2204 7062 2976
rect 7050 2196 7052 2204
rect 7060 2196 7062 2204
rect 7050 2194 7062 2196
rect 7082 2924 7094 2926
rect 7082 2916 7084 2924
rect 7092 2916 7094 2924
rect 7050 1884 7062 1886
rect 7050 1876 7052 1884
rect 7060 1876 7062 1884
rect 7050 1124 7062 1876
rect 7050 1116 7052 1124
rect 7060 1116 7062 1124
rect 7050 1114 7062 1116
rect 7082 744 7094 2916
rect 7178 2844 7190 2846
rect 7178 2836 7180 2844
rect 7188 2836 7190 2844
rect 7146 2724 7158 2726
rect 7146 2716 7148 2724
rect 7156 2716 7158 2724
rect 7114 2124 7126 2126
rect 7114 2116 7116 2124
rect 7124 2116 7126 2124
rect 7114 2004 7126 2116
rect 7114 1996 7116 2004
rect 7124 1996 7126 2004
rect 7114 1994 7126 1996
rect 7114 1884 7126 1886
rect 7114 1876 7116 1884
rect 7124 1876 7126 1884
rect 7114 1484 7126 1876
rect 7146 1784 7158 2716
rect 7178 2224 7190 2836
rect 7178 2216 7180 2224
rect 7188 2216 7190 2224
rect 7178 2214 7190 2216
rect 7210 2384 7222 2386
rect 7210 2376 7212 2384
rect 7220 2376 7222 2384
rect 7146 1776 7148 1784
rect 7156 1776 7158 1784
rect 7146 1774 7158 1776
rect 7178 2044 7190 2046
rect 7178 2036 7180 2044
rect 7188 2036 7190 2044
rect 7178 1784 7190 2036
rect 7178 1776 7180 1784
rect 7188 1776 7190 1784
rect 7114 1476 7116 1484
rect 7124 1476 7126 1484
rect 7114 1474 7126 1476
rect 7146 1744 7158 1746
rect 7146 1736 7148 1744
rect 7156 1736 7158 1744
rect 7146 1424 7158 1736
rect 7178 1644 7190 1776
rect 7178 1636 7180 1644
rect 7188 1636 7190 1644
rect 7178 1634 7190 1636
rect 7146 1416 7148 1424
rect 7156 1416 7158 1424
rect 7146 1414 7158 1416
rect 7178 1584 7190 1586
rect 7178 1576 7180 1584
rect 7188 1576 7190 1584
rect 7082 736 7084 744
rect 7092 736 7094 744
rect 7082 734 7094 736
rect 7114 964 7126 966
rect 7114 956 7116 964
rect 7124 956 7126 964
rect 7114 544 7126 956
rect 7114 536 7116 544
rect 7124 536 7126 544
rect 7114 534 7126 536
rect 7178 444 7190 1576
rect 7210 684 7222 2376
rect 7242 1544 7254 3756
rect 7274 3244 7286 4596
rect 7274 3236 7276 3244
rect 7284 3236 7286 3244
rect 7274 3234 7286 3236
rect 7242 1536 7244 1544
rect 7252 1536 7254 1544
rect 7242 1534 7254 1536
rect 7274 2524 7286 2526
rect 7274 2516 7276 2524
rect 7284 2516 7286 2524
rect 7242 1504 7254 1506
rect 7242 1496 7244 1504
rect 7252 1496 7254 1504
rect 7242 924 7254 1496
rect 7242 916 7244 924
rect 7252 916 7254 924
rect 7242 914 7254 916
rect 7274 904 7286 2516
rect 7306 1904 7318 5036
rect 7338 3784 7350 3786
rect 7338 3776 7340 3784
rect 7348 3776 7350 3784
rect 7338 2764 7350 3776
rect 7338 2756 7340 2764
rect 7348 2756 7350 2764
rect 7338 2754 7350 2756
rect 7306 1896 7308 1904
rect 7316 1896 7318 1904
rect 7306 1894 7318 1896
rect 7338 2704 7350 2706
rect 7338 2696 7340 2704
rect 7348 2696 7350 2704
rect 7306 1864 7318 1866
rect 7306 1856 7308 1864
rect 7316 1856 7318 1864
rect 7306 1564 7318 1856
rect 7338 1844 7350 2696
rect 7370 2364 7382 5076
rect 7402 3324 7414 3326
rect 7402 3316 7404 3324
rect 7412 3316 7414 3324
rect 7402 2824 7414 3316
rect 7402 2816 7404 2824
rect 7412 2816 7414 2824
rect 7402 2814 7414 2816
rect 7370 2356 7372 2364
rect 7380 2356 7382 2364
rect 7370 2354 7382 2356
rect 7338 1836 7340 1844
rect 7348 1836 7350 1844
rect 7338 1834 7350 1836
rect 7370 2304 7382 2306
rect 7370 2296 7372 2304
rect 7380 2296 7382 2304
rect 7306 1556 7308 1564
rect 7316 1556 7318 1564
rect 7306 1554 7318 1556
rect 7338 1764 7350 1766
rect 7338 1756 7340 1764
rect 7348 1756 7350 1764
rect 7306 1084 7318 1086
rect 7306 1076 7308 1084
rect 7316 1076 7318 1084
rect 7306 1044 7318 1076
rect 7306 1036 7308 1044
rect 7316 1036 7318 1044
rect 7306 1034 7318 1036
rect 7274 896 7276 904
rect 7284 896 7286 904
rect 7274 894 7286 896
rect 7306 1004 7318 1006
rect 7306 996 7308 1004
rect 7316 996 7318 1004
rect 7210 676 7212 684
rect 7220 676 7222 684
rect 7210 674 7222 676
rect 7306 644 7318 996
rect 7338 664 7350 1756
rect 7370 1024 7382 2296
rect 7370 1016 7372 1024
rect 7380 1016 7382 1024
rect 7370 1014 7382 1016
rect 7402 2244 7414 2246
rect 7402 2236 7404 2244
rect 7412 2236 7414 2244
rect 7338 656 7340 664
rect 7348 656 7350 664
rect 7338 654 7350 656
rect 7370 984 7382 986
rect 7370 976 7372 984
rect 7380 976 7382 984
rect 7306 636 7308 644
rect 7316 636 7318 644
rect 7306 634 7318 636
rect 7178 436 7180 444
rect 7188 436 7190 444
rect 7178 434 7190 436
rect 7370 304 7382 976
rect 7402 324 7414 2236
rect 7402 316 7404 324
rect 7412 316 7414 324
rect 7402 314 7414 316
rect 7370 296 7372 304
rect 7380 296 7382 304
rect 7370 294 7382 296
rect 7018 136 7020 144
rect 7028 136 7030 144
rect 7018 134 7030 136
rect 6634 96 6636 104
rect 6644 96 6646 104
rect 6634 94 6646 96
use INVX1  _2438_
timestamp 1596033377
transform 1 0 8 0 -1 210
box -4 -6 36 206
use NOR2X1  _2447_
timestamp 1596033377
transform 1 0 40 0 -1 210
box -4 -6 52 206
use NAND2X1  _2437_
timestamp 1596033377
transform 1 0 88 0 -1 210
box -4 -6 52 206
use INVX1  _2436_
timestamp 1596033377
transform -1 0 168 0 -1 210
box -4 -6 36 206
use NAND2X1  _2439_
timestamp 1596033377
transform 1 0 168 0 -1 210
box -4 -6 52 206
use XNOR2X1  _2441_
timestamp 1596033377
transform 1 0 8 0 1 210
box -4 -6 116 206
use OAI21X1  _2448_
timestamp 1596033377
transform 1 0 120 0 1 210
box -4 -6 68 206
use NAND2X1  _2440_
timestamp 1596033377
transform 1 0 184 0 1 210
box -4 -6 52 206
use NOR2X1  _2442_
timestamp 1596033377
transform -1 0 344 0 1 210
box -4 -6 52 206
use AOI21X1  _2443_
timestamp 1596033377
transform 1 0 232 0 1 210
box -4 -6 68 206
use NAND2X1  _2435_
timestamp 1596033377
transform -1 0 328 0 -1 210
box -4 -6 52 206
use AND2X2  _2446_
timestamp 1596033377
transform -1 0 280 0 -1 210
box -4 -6 68 206
use INVX1  _2799_
timestamp 1596033377
transform -1 0 408 0 1 210
box -4 -6 36 206
use INVX1  _2797_
timestamp 1596033377
transform 1 0 344 0 1 210
box -4 -6 36 206
use NAND2X1  _2803_
timestamp 1596033377
transform -1 0 408 0 -1 210
box -4 -6 52 206
use INVX1  _2434_
timestamp 1596033377
transform -1 0 360 0 -1 210
box -4 -6 36 206
use OAI22X1  _2798_
timestamp 1596033377
transform -1 0 488 0 1 210
box -4 -6 84 206
use NOR2X1  _2805_
timestamp 1596033377
transform 1 0 408 0 -1 210
box -4 -6 52 206
use OAI21X1  _2806_
timestamp 1596033377
transform -1 0 520 0 -1 210
box -4 -6 68 206
use BUFX2  _2096_
timestamp 1596033377
transform 1 0 520 0 -1 210
box -4 -6 52 206
use INVX1  _2790_
timestamp 1596033377
transform 1 0 568 0 -1 210
box -4 -6 36 206
use NAND2X1  _2791_
timestamp 1596033377
transform 1 0 600 0 -1 210
box -4 -6 52 206
use INVX1  _2796_
timestamp 1596033377
transform -1 0 520 0 1 210
box -4 -6 36 206
use OAI22X1  _2801_
timestamp 1596033377
transform 1 0 520 0 1 210
box -4 -6 84 206
use NAND2X1  _2804_
timestamp 1596033377
transform 1 0 600 0 1 210
box -4 -6 52 206
use NOR2X1  _2792_
timestamp 1596033377
transform -1 0 696 0 -1 210
box -4 -6 52 206
use BUFX2  _2097_
timestamp 1596033377
transform -1 0 744 0 -1 210
box -4 -6 52 206
use NOR2X1  _2903_
timestamp 1596033377
transform 1 0 744 0 -1 210
box -4 -6 52 206
use INVX1  _2902_
timestamp 1596033377
transform 1 0 792 0 -1 210
box -4 -6 36 206
use INVX1  _2800_
timestamp 1596033377
transform -1 0 680 0 1 210
box -4 -6 36 206
use NOR2X1  _2802_
timestamp 1596033377
transform -1 0 728 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert168
timestamp 1596033377
transform -1 0 776 0 1 210
box -4 -6 52 206
use INVX1  _2793_
timestamp 1596033377
transform 1 0 776 0 1 210
box -4 -6 36 206
use OAI21X1  _2840_
timestamp 1596033377
transform -1 0 872 0 1 210
box -4 -6 68 206
use NAND2X1  _2906_
timestamp 1596033377
transform -1 0 872 0 -1 210
box -4 -6 52 206
use AOI21X1  _2907_
timestamp 1596033377
transform -1 0 936 0 -1 210
box -4 -6 68 206
use NAND2X1  _2905_
timestamp 1596033377
transform 1 0 936 0 -1 210
box -4 -6 52 206
use INVX1  _2904_
timestamp 1596033377
transform -1 0 1016 0 -1 210
box -4 -6 36 206
use NOR2X1  _2794_
timestamp 1596033377
transform -1 0 920 0 1 210
box -4 -6 52 206
use OAI21X1  _2795_
timestamp 1596033377
transform -1 0 984 0 1 210
box -4 -6 68 206
use NOR2X1  _2841_
timestamp 1596033377
transform -1 0 1032 0 1 210
box -4 -6 52 206
use XNOR2X1  _2463_
timestamp 1596033377
transform 1 0 1016 0 -1 210
box -4 -6 116 206
use XOR2X1  _2460_
timestamp 1596033377
transform -1 0 1240 0 -1 210
box -4 -6 116 206
use BUFX2  BUFX2_insert171
timestamp 1596033377
transform 1 0 1032 0 1 210
box -4 -6 52 206
use AOI21X1  _2807_
timestamp 1596033377
transform -1 0 1144 0 1 210
box -4 -6 68 206
use OAI21X1  _2842_
timestamp 1596033377
transform -1 0 1208 0 1 210
box -4 -6 68 206
use INVX1  _2838_
timestamp 1596033377
transform 1 0 1208 0 1 210
box -4 -6 36 206
use NAND2X1  _2485_
timestamp 1596033377
transform 1 0 1240 0 -1 210
box -4 -6 52 206
use INVX1  _2466_
timestamp 1596033377
transform -1 0 1320 0 -1 210
box -4 -6 36 206
use NAND2X1  _2467_
timestamp 1596033377
transform -1 0 1368 0 -1 210
box -4 -6 52 206
use NAND2X1  _2464_
timestamp 1596033377
transform 1 0 1240 0 1 210
box -4 -6 52 206
use NOR2X1  _2473_
timestamp 1596033377
transform 1 0 1288 0 1 210
box -4 -6 52 206
use NOR3X1  _2843_
timestamp 1596033377
transform -1 0 1464 0 1 210
box -4 -6 132 206
use FILL  SFILL13680x100
timestamp 1596033377
transform -1 0 1384 0 -1 210
box -4 -6 20 206
use FILL  SFILL13840x100
timestamp 1596033377
transform -1 0 1400 0 -1 210
box -4 -6 20 206
use FILL  SFILL14000x100
timestamp 1596033377
transform -1 0 1416 0 -1 210
box -4 -6 20 206
use FILL  SFILL14960x2100
timestamp 1596033377
transform 1 0 1496 0 1 210
box -4 -6 20 206
use FILL  SFILL14800x2100
timestamp 1596033377
transform 1 0 1480 0 1 210
box -4 -6 20 206
use FILL  SFILL14640x2100
timestamp 1596033377
transform 1 0 1464 0 1 210
box -4 -6 20 206
use FILL  SFILL14160x100
timestamp 1596033377
transform -1 0 1432 0 -1 210
box -4 -6 20 206
use FILL  SFILL15120x2100
timestamp 1596033377
transform 1 0 1512 0 1 210
box -4 -6 20 206
use NAND2X1  _2470_
timestamp 1596033377
transform 1 0 1592 0 1 210
box -4 -6 52 206
use OAI21X1  _2825_
timestamp 1596033377
transform 1 0 1528 0 1 210
box -4 -6 68 206
use AOI21X1  _2820_
timestamp 1596033377
transform 1 0 1576 0 -1 210
box -4 -6 68 206
use INVX1  _2818_
timestamp 1596033377
transform 1 0 1544 0 -1 210
box -4 -6 36 206
use XNOR2X1  _2484_
timestamp 1596033377
transform -1 0 1544 0 -1 210
box -4 -6 116 206
use NAND3X1  _2821_
timestamp 1596033377
transform -1 0 1704 0 -1 210
box -4 -6 68 206
use NOR2X1  _2819_
timestamp 1596033377
transform 1 0 1704 0 -1 210
box -4 -6 52 206
use INVX1  _2462_
timestamp 1596033377
transform 1 0 1752 0 -1 210
box -4 -6 36 206
use INVX1  _2815_
timestamp 1596033377
transform -1 0 1816 0 -1 210
box -4 -6 36 206
use INVX1  _2468_
timestamp 1596033377
transform -1 0 1672 0 1 210
box -4 -6 36 206
use NAND2X1  _2469_
timestamp 1596033377
transform -1 0 1720 0 1 210
box -4 -6 52 206
use OAI21X1  _2472_
timestamp 1596033377
transform -1 0 1784 0 1 210
box -4 -6 68 206
use OAI21X1  _2465_
timestamp 1596033377
transform 1 0 1784 0 1 210
box -4 -6 68 206
use NOR2X1  _2823_
timestamp 1596033377
transform 1 0 1816 0 -1 210
box -4 -6 52 206
use AOI22X1  _2817_
timestamp 1596033377
transform 1 0 1864 0 -1 210
box -4 -6 84 206
use INVX1  _2816_
timestamp 1596033377
transform -1 0 1976 0 -1 210
box -4 -6 36 206
use AOI22X1  _2606_
timestamp 1596033377
transform 1 0 1976 0 -1 210
box -4 -6 84 206
use AOI22X1  _2824_
timestamp 1596033377
transform -1 0 1928 0 1 210
box -4 -6 84 206
use NAND2X1  _2822_
timestamp 1596033377
transform -1 0 1976 0 1 210
box -4 -6 52 206
use NOR2X1  _2814_
timestamp 1596033377
transform 1 0 1976 0 1 210
box -4 -6 52 206
use INVX1  _2605_
timestamp 1596033377
transform -1 0 2088 0 -1 210
box -4 -6 36 206
use OAI22X1  _2632_
timestamp 1596033377
transform -1 0 2168 0 -1 210
box -4 -6 84 206
use INVX1  _2604_
timestamp 1596033377
transform -1 0 2200 0 -1 210
box -4 -6 36 206
use BUFX2  _2106_
timestamp 1596033377
transform -1 0 2248 0 -1 210
box -4 -6 52 206
use XNOR2X1  _2471_
timestamp 1596033377
transform -1 0 2136 0 1 210
box -4 -6 116 206
use INVX1  _3098_
timestamp 1596033377
transform 1 0 2136 0 1 210
box -4 -6 36 206
use BUFX2  BUFX2_insert287
timestamp 1596033377
transform -1 0 2216 0 1 210
box -4 -6 52 206
use INVX1  _2700_
timestamp 1596033377
transform 1 0 2248 0 -1 210
box -4 -6 36 206
use NAND2X1  _2701_
timestamp 1596033377
transform 1 0 2280 0 -1 210
box -4 -6 52 206
use OAI22X1  _2722_
timestamp 1596033377
transform -1 0 2408 0 -1 210
box -4 -6 84 206
use INVX1  _2698_
timestamp 1596033377
transform 1 0 2408 0 -1 210
box -4 -6 36 206
use NAND2X1  _2607_
timestamp 1596033377
transform -1 0 2264 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert268
timestamp 1596033377
transform -1 0 2312 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert157
timestamp 1596033377
transform -1 0 2360 0 1 210
box -4 -6 52 206
use OAI21X1  _2633_
timestamp 1596033377
transform -1 0 2424 0 1 210
box -4 -6 68 206
use NAND2X1  _2699_
timestamp 1596033377
transform -1 0 2488 0 -1 210
box -4 -6 52 206
use BUFX2  _2107_
timestamp 1596033377
transform -1 0 2536 0 -1 210
box -4 -6 52 206
use BUFX2  _2109_
timestamp 1596033377
transform -1 0 2584 0 -1 210
box -4 -6 52 206
use OAI22X1  _2813_
timestamp 1596033377
transform 1 0 2584 0 -1 210
box -4 -6 84 206
use BUFX2  BUFX2_insert55
timestamp 1596033377
transform -1 0 2472 0 1 210
box -4 -6 52 206
use NAND3X1  _2702_
timestamp 1596033377
transform 1 0 2472 0 1 210
box -4 -6 68 206
use INVX1  _2601_
timestamp 1596033377
transform 1 0 2536 0 1 210
box -4 -6 36 206
use AOI22X1  _2603_
timestamp 1596033377
transform 1 0 2568 0 1 210
box -4 -6 84 206
use INVX1  _2811_
timestamp 1596033377
transform -1 0 2696 0 -1 210
box -4 -6 36 206
use INVX1  _2812_
timestamp 1596033377
transform -1 0 2728 0 -1 210
box -4 -6 36 206
use INVX1  _2689_
timestamp 1596033377
transform 1 0 2728 0 -1 210
box -4 -6 36 206
use NOR2X1  _2726_
timestamp 1596033377
transform 1 0 2760 0 -1 210
box -4 -6 52 206
use AOI22X1  _2690_
timestamp 1596033377
transform -1 0 2888 0 -1 210
box -4 -6 84 206
use INVX1  _2602_
timestamp 1596033377
transform -1 0 2680 0 1 210
box -4 -6 36 206
use INVX1  _2696_
timestamp 1596033377
transform 1 0 2680 0 1 210
box -4 -6 36 206
use AOI22X1  _2697_
timestamp 1596033377
transform -1 0 2792 0 1 210
box -4 -6 84 206
use INVX1  _2695_
timestamp 1596033377
transform 1 0 2792 0 1 210
box -4 -6 36 206
use OAI21X1  _2723_
timestamp 1596033377
transform 1 0 2824 0 1 210
box -4 -6 68 206
use FILL  SFILL29520x2100
timestamp 1596033377
transform 1 0 2952 0 1 210
box -4 -6 20 206
use FILL  SFILL29520x100
timestamp 1596033377
transform -1 0 2968 0 -1 210
box -4 -6 20 206
use FILL  SFILL29360x100
timestamp 1596033377
transform -1 0 2952 0 -1 210
box -4 -6 20 206
use FILL  SFILL29200x100
timestamp 1596033377
transform -1 0 2936 0 -1 210
box -4 -6 20 206
use OAI21X1  _2728_
timestamp 1596033377
transform 1 0 2888 0 1 210
box -4 -6 68 206
use INVX1  _2688_
timestamp 1596033377
transform -1 0 2920 0 -1 210
box -4 -6 36 206
use FILL  SFILL30000x2100
timestamp 1596033377
transform 1 0 3000 0 1 210
box -4 -6 20 206
use FILL  SFILL29840x2100
timestamp 1596033377
transform 1 0 2984 0 1 210
box -4 -6 20 206
use FILL  SFILL29680x2100
timestamp 1596033377
transform 1 0 2968 0 1 210
box -4 -6 20 206
use FILL  SFILL29680x100
timestamp 1596033377
transform -1 0 2984 0 -1 210
box -4 -6 20 206
use AOI21X1  _2727_
timestamp 1596033377
transform 1 0 2984 0 -1 210
box -4 -6 68 206
use BUFX2  _2108_
timestamp 1596033377
transform 1 0 3048 0 -1 210
box -4 -6 52 206
use BUFX2  _2088_
timestamp 1596033377
transform -1 0 3144 0 -1 210
box -4 -6 52 206
use BUFX2  _2092_
timestamp 1596033377
transform 1 0 3144 0 -1 210
box -4 -6 52 206
use BUFX2  _2091_
timestamp 1596033377
transform -1 0 3240 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert54
timestamp 1596033377
transform -1 0 3064 0 1 210
box -4 -6 52 206
use NAND2X1  _2694_
timestamp 1596033377
transform 1 0 3064 0 1 210
box -4 -6 52 206
use NOR2X1  _2724_
timestamp 1596033377
transform -1 0 3160 0 1 210
box -4 -6 52 206
use INVX1  _2691_
timestamp 1596033377
transform 1 0 3160 0 1 210
box -4 -6 36 206
use NAND2X1  _2725_
timestamp 1596033377
transform -1 0 3240 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3636_
timestamp 1596033377
transform -1 0 3432 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert267
timestamp 1596033377
transform 1 0 3240 0 1 210
box -4 -6 52 206
use AOI22X1  _2693_
timestamp 1596033377
transform 1 0 3288 0 1 210
box -4 -6 84 206
use INVX1  _2692_
timestamp 1596033377
transform 1 0 3368 0 1 210
box -4 -6 36 206
use DFFPOSX1  _3637_
timestamp 1596033377
transform -1 0 3592 0 1 210
box -4 -6 196 206
use DFFPOSX1  _3421_
timestamp 1596033377
transform 1 0 3432 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _3419_
timestamp 1596033377
transform 1 0 3592 0 1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert131
timestamp 1596033377
transform 1 0 3624 0 -1 210
box -4 -6 52 206
use BUFX2  _2112_
timestamp 1596033377
transform 1 0 3672 0 -1 210
box -4 -6 52 206
use NAND2X1  _3598_
timestamp 1596033377
transform 1 0 3720 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3630_
timestamp 1596033377
transform 1 0 3768 0 -1 210
box -4 -6 196 206
use AOI21X1  _3600_
timestamp 1596033377
transform 1 0 3784 0 1 210
box -4 -6 68 206
use NAND2X1  _3607_
timestamp 1596033377
transform 1 0 3960 0 -1 210
box -4 -6 52 206
use AOI21X1  _3609_
timestamp 1596033377
transform -1 0 4072 0 -1 210
box -4 -6 68 206
use NAND2X1  _3599_
timestamp 1596033377
transform 1 0 3848 0 1 210
box -4 -6 52 206
use INVX1  _3381_
timestamp 1596033377
transform 1 0 3896 0 1 210
box -4 -6 36 206
use AOI21X1  _3603_
timestamp 1596033377
transform -1 0 3992 0 1 210
box -4 -6 68 206
use NAND2X1  _3602_
timestamp 1596033377
transform -1 0 4040 0 1 210
box -4 -6 52 206
use NAND2X1  _3595_
timestamp 1596033377
transform 1 0 4072 0 -1 210
box -4 -6 52 206
use AOI21X1  _3597_
timestamp 1596033377
transform 1 0 4120 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _3626_
timestamp 1596033377
transform 1 0 4184 0 -1 210
box -4 -6 196 206
use NAND2X1  _3601_
timestamp 1596033377
transform -1 0 4088 0 1 210
box -4 -6 52 206
use INVX1  _3437_
timestamp 1596033377
transform 1 0 4088 0 1 210
box -4 -6 36 206
use NAND2X1  _3596_
timestamp 1596033377
transform -1 0 4168 0 1 210
box -4 -6 52 206
use NAND2X1  _3608_
timestamp 1596033377
transform -1 0 4216 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3635_
timestamp 1596033377
transform -1 0 4408 0 1 210
box -4 -6 196 206
use AOI21X1  _3606_
timestamp 1596033377
transform -1 0 4440 0 -1 210
box -4 -6 68 206
use FILL  SFILL44080x2100
timestamp 1596033377
transform 1 0 4408 0 1 210
box -4 -6 20 206
use FILL  SFILL44560x2100
timestamp 1596033377
transform 1 0 4456 0 1 210
box -4 -6 20 206
use FILL  SFILL44400x2100
timestamp 1596033377
transform 1 0 4440 0 1 210
box -4 -6 20 206
use FILL  SFILL44240x2100
timestamp 1596033377
transform 1 0 4424 0 1 210
box -4 -6 20 206
use FILL  SFILL44880x100
timestamp 1596033377
transform -1 0 4504 0 -1 210
box -4 -6 20 206
use FILL  SFILL44720x100
timestamp 1596033377
transform -1 0 4488 0 -1 210
box -4 -6 20 206
use FILL  SFILL44560x100
timestamp 1596033377
transform -1 0 4472 0 -1 210
box -4 -6 20 206
use FILL  SFILL44400x100
timestamp 1596033377
transform -1 0 4456 0 -1 210
box -4 -6 20 206
use BUFX2  BUFX2_insert134
timestamp 1596033377
transform 1 0 4504 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert132
timestamp 1596033377
transform 1 0 4600 0 -1 210
box -4 -6 52 206
use NAND2X1  _3604_
timestamp 1596033377
transform 1 0 4552 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _3627_
timestamp 1596033377
transform -1 0 4664 0 1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert133
timestamp 1596033377
transform 1 0 4648 0 -1 210
box -4 -6 52 206
use NAND2X1  _3572_
timestamp 1596033377
transform 1 0 4696 0 -1 210
box -4 -6 52 206
use NAND2X1  _3578_
timestamp 1596033377
transform 1 0 4744 0 -1 210
box -4 -6 52 206
use NAND2X1  _3581_
timestamp 1596033377
transform 1 0 4792 0 -1 210
box -4 -6 52 206
use NAND2X1  _3614_
timestamp 1596033377
transform 1 0 4664 0 1 210
box -4 -6 52 206
use INVX1  _3458_
timestamp 1596033377
transform -1 0 4744 0 1 210
box -4 -6 36 206
use AOI21X1  _3615_
timestamp 1596033377
transform 1 0 4744 0 1 210
box -4 -6 68 206
use INVX1  _3472_
timestamp 1596033377
transform -1 0 4840 0 1 210
box -4 -6 36 206
use DFFPOSX1  _3646_
timestamp 1596033377
transform -1 0 5032 0 -1 210
box -4 -6 196 206
use INVX1  _3428_
timestamp 1596033377
transform 1 0 4840 0 1 210
box -4 -6 36 206
use NAND2X1  _3605_
timestamp 1596033377
transform 1 0 4872 0 1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert124
timestamp 1596033377
transform -1 0 4968 0 1 210
box -4 -6 52 206
use INVX1  _3500_
timestamp 1596033377
transform -1 0 5000 0 1 210
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert24
timestamp 1596033377
transform -1 0 5144 0 1 210
box -4 -6 148 206
use NAND2X1  _3583_
timestamp 1596033377
transform 1 0 5032 0 -1 210
box -4 -6 52 206
use NAND2X1  _3566_
timestamp 1596033377
transform 1 0 5080 0 -1 210
box -4 -6 52 206
use NAND2X1  _3586_
timestamp 1596033377
transform 1 0 5128 0 -1 210
box -4 -6 52 206
use NAND2X1  _3589_
timestamp 1596033377
transform 1 0 5176 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_insert19
timestamp 1596033377
transform -1 0 5192 0 1 210
box -4 -6 52 206
use INVX8  _3564_
timestamp 1596033377
transform 1 0 5192 0 1 210
box -4 -6 84 206
use AOI21X1  _3582_
timestamp 1596033377
transform 1 0 5224 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _3643_
timestamp 1596033377
transform 1 0 5288 0 -1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert126
timestamp 1596033377
transform 1 0 5272 0 1 210
box -4 -6 52 206
use AOI21X1  _3573_
timestamp 1596033377
transform -1 0 5384 0 1 210
box -4 -6 68 206
use BUFX2  BUFX2_insert18
timestamp 1596033377
transform 1 0 5384 0 1 210
box -4 -6 52 206
use DFFPOSX1  _3639_
timestamp 1596033377
transform 1 0 5480 0 -1 210
box -4 -6 196 206
use NAND2X1  _3571_
timestamp 1596033377
transform -1 0 5480 0 1 210
box -4 -6 52 206
use INVX8  _3905_
timestamp 1596033377
transform 1 0 5480 0 1 210
box -4 -6 84 206
use NAND2X1  _3565_
timestamp 1596033377
transform 1 0 5560 0 1 210
box -4 -6 52 206
use AOI21X1  _3567_
timestamp 1596033377
transform 1 0 5608 0 1 210
box -4 -6 68 206
use AOI21X1  _3585_
timestamp 1596033377
transform -1 0 5736 0 -1 210
box -4 -6 68 206
use DFFPOSX1  _3638_
timestamp 1596033377
transform 1 0 5736 0 -1 210
box -4 -6 196 206
use AOI21X1  _3588_
timestamp 1596033377
transform -1 0 5736 0 1 210
box -4 -6 68 206
use NAND2X1  _3580_
timestamp 1596033377
transform -1 0 5784 0 1 210
box -4 -6 52 206
use NAND2X1  _3587_
timestamp 1596033377
transform -1 0 5832 0 1 210
box -4 -6 52 206
use INVX8  _4085_
timestamp 1596033377
transform 1 0 5880 0 1 210
box -4 -6 84 206
use NAND2X1  _3584_
timestamp 1596033377
transform -1 0 5880 0 1 210
box -4 -6 52 206
use FILL  SFILL59920x2100
timestamp 1596033377
transform 1 0 5992 0 1 210
box -4 -6 20 206
use FILL  SFILL59760x2100
timestamp 1596033377
transform 1 0 5976 0 1 210
box -4 -6 20 206
use FILL  SFILL59600x2100
timestamp 1596033377
transform 1 0 5960 0 1 210
box -4 -6 20 206
use FILL  SFILL59760x100
timestamp 1596033377
transform -1 0 5992 0 -1 210
box -4 -6 20 206
use FILL  SFILL59600x100
timestamp 1596033377
transform -1 0 5976 0 -1 210
box -4 -6 20 206
use FILL  SFILL59440x100
timestamp 1596033377
transform -1 0 5960 0 -1 210
box -4 -6 20 206
use FILL  SFILL59280x100
timestamp 1596033377
transform -1 0 5944 0 -1 210
box -4 -6 20 206
use AOI21X1  _3668_
timestamp 1596033377
transform 1 0 5992 0 -1 210
box -4 -6 68 206
use FILL  SFILL60080x2100
timestamp 1596033377
transform 1 0 6008 0 1 210
box -4 -6 20 206
use NOR2X1  _3667_
timestamp 1596033377
transform -1 0 6104 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _4397_
timestamp 1596033377
transform 1 0 6104 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _3644_
timestamp 1596033377
transform 1 0 6024 0 1 210
box -4 -6 196 206
use BUFX2  BUFX2_insert86
timestamp 1596033377
transform 1 0 6216 0 1 210
box -4 -6 52 206
use DFFPOSX1  _4381_
timestamp 1596033377
transform 1 0 6296 0 -1 210
box -4 -6 196 206
use OAI21X1  _3851_
timestamp 1596033377
transform 1 0 6264 0 1 210
box -4 -6 68 206
use NAND2X1  _3850_
timestamp 1596033377
transform -1 0 6376 0 1 210
box -4 -6 52 206
use DFFPOSX1  _4301_
timestamp 1596033377
transform 1 0 6376 0 1 210
box -4 -6 196 206
use DFFPOSX1  _4330_
timestamp 1596033377
transform -1 0 6680 0 -1 210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert27
timestamp 1596033377
transform -1 0 6712 0 1 210
box -4 -6 148 206
use DFFPOSX1  _4371_
timestamp 1596033377
transform -1 0 6872 0 -1 210
box -4 -6 196 206
use OAI21X1  _3784_
timestamp 1596033377
transform 1 0 6712 0 1 210
box -4 -6 68 206
use DFFPOSX1  _4349_
timestamp 1596033377
transform 1 0 6776 0 1 210
box -4 -6 196 206
use DFFPOSX1  _4405_
timestamp 1596033377
transform 1 0 6872 0 -1 210
box -4 -6 196 206
use OAI21X1  _3719_
timestamp 1596033377
transform -1 0 7032 0 1 210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert33
timestamp 1596033377
transform -1 0 7208 0 -1 210
box -4 -6 148 206
use CLKBUF1  CLKBUF1_insert26
timestamp 1596033377
transform -1 0 7352 0 -1 210
box -4 -6 148 206
use CLKBUF1  CLKBUF1_insert34
timestamp 1596033377
transform 1 0 7032 0 1 210
box -4 -6 148 206
use DFFPOSX1  _4382_
timestamp 1596033377
transform 1 0 7176 0 1 210
box -4 -6 196 206
use FILL  FILL70960x100
timestamp 1596033377
transform -1 0 7368 0 -1 210
box -4 -6 20 206
use FILL  FILL71120x100
timestamp 1596033377
transform -1 0 7384 0 -1 210
box -4 -6 20 206
use FILL  FILL71280x100
timestamp 1596033377
transform -1 0 7400 0 -1 210
box -4 -6 20 206
use FILL  FILL71120x2100
timestamp 1596033377
transform 1 0 7368 0 1 210
box -4 -6 20 206
use FILL  FILL71280x2100
timestamp 1596033377
transform 1 0 7384 0 1 210
box -4 -6 20 206
use NOR2X1  _2450_
timestamp 1596033377
transform -1 0 56 0 -1 610
box -4 -6 52 206
use INVX1  _2449_
timestamp 1596033377
transform -1 0 88 0 -1 610
box -4 -6 36 206
use XNOR2X1  _2444_
timestamp 1596033377
transform 1 0 88 0 -1 610
box -4 -6 116 206
use OAI21X1  _2459_
timestamp 1596033377
transform -1 0 264 0 -1 610
box -4 -6 68 206
use AOI21X1  _2458_
timestamp 1596033377
transform 1 0 264 0 -1 610
box -4 -6 68 206
use NOR2X1  _2457_
timestamp 1596033377
transform -1 0 376 0 -1 610
box -4 -6 52 206
use NAND2X1  _2456_
timestamp 1596033377
transform -1 0 424 0 -1 610
box -4 -6 52 206
use INVX1  _2455_
timestamp 1596033377
transform -1 0 456 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert96
timestamp 1596033377
transform -1 0 504 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert247
timestamp 1596033377
transform -1 0 552 0 -1 610
box -4 -6 52 206
use AOI21X1  _2625_
timestamp 1596033377
transform -1 0 616 0 -1 610
box -4 -6 68 206
use NAND2X1  _2620_
timestamp 1596033377
transform 1 0 616 0 -1 610
box -4 -6 52 206
use NOR2X1  _2624_
timestamp 1596033377
transform -1 0 712 0 -1 610
box -4 -6 52 206
use NAND2X1  _2617_
timestamp 1596033377
transform -1 0 760 0 -1 610
box -4 -6 52 206
use INVX1  _2616_
timestamp 1596033377
transform -1 0 792 0 -1 610
box -4 -6 36 206
use OAI22X1  _2621_
timestamp 1596033377
transform 1 0 792 0 -1 610
box -4 -6 84 206
use NAND2X1  _2619_
timestamp 1596033377
transform -1 0 920 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert297
timestamp 1596033377
transform -1 0 968 0 -1 610
box -4 -6 52 206
use INVX1  _2618_
timestamp 1596033377
transform -1 0 1000 0 -1 610
box -4 -6 36 206
use AOI21X1  _2493_
timestamp 1596033377
transform -1 0 1064 0 -1 610
box -4 -6 68 206
use XNOR2X1  _2461_
timestamp 1596033377
transform 1 0 1064 0 -1 610
box -4 -6 116 206
use INVX1  _2839_
timestamp 1596033377
transform 1 0 1176 0 -1 610
box -4 -6 36 206
use NOR2X1  _2487_
timestamp 1596033377
transform 1 0 1208 0 -1 610
box -4 -6 52 206
use OAI21X1  _2492_
timestamp 1596033377
transform 1 0 1256 0 -1 610
box -4 -6 68 206
use AOI22X1  _2474_
timestamp 1596033377
transform -1 0 1400 0 -1 610
box -4 -6 84 206
use FILL  SFILL14000x4100
timestamp 1596033377
transform -1 0 1416 0 -1 610
box -4 -6 20 206
use OAI21X1  _2488_
timestamp 1596033377
transform -1 0 1528 0 -1 610
box -4 -6 68 206
use XOR2X1  _2479_
timestamp 1596033377
transform 1 0 1528 0 -1 610
box -4 -6 116 206
use FILL  SFILL14160x4100
timestamp 1596033377
transform -1 0 1432 0 -1 610
box -4 -6 20 206
use FILL  SFILL14320x4100
timestamp 1596033377
transform -1 0 1448 0 -1 610
box -4 -6 20 206
use FILL  SFILL14480x4100
timestamp 1596033377
transform -1 0 1464 0 -1 610
box -4 -6 20 206
use AOI21X1  _2491_
timestamp 1596033377
transform -1 0 1704 0 -1 610
box -4 -6 68 206
use NOR2X1  _2490_
timestamp 1596033377
transform 1 0 1704 0 -1 610
box -4 -6 52 206
use INVX1  _2489_
timestamp 1596033377
transform -1 0 1784 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert82
timestamp 1596033377
transform -1 0 1832 0 -1 610
box -4 -6 52 206
use INVX1  _2808_
timestamp 1596033377
transform 1 0 1832 0 -1 610
box -4 -6 36 206
use OAI22X1  _2810_
timestamp 1596033377
transform 1 0 1864 0 -1 610
box -4 -6 84 206
use INVX1  _2595_
timestamp 1596033377
transform 1 0 1944 0 -1 610
box -4 -6 36 206
use AOI22X1  _2596_
timestamp 1596033377
transform -1 0 2056 0 -1 610
box -4 -6 84 206
use NOR2X1  _2631_
timestamp 1596033377
transform -1 0 2104 0 -1 610
box -4 -6 52 206
use OAI22X1  _2634_
timestamp 1596033377
transform 1 0 2104 0 -1 610
box -4 -6 84 206
use NOR2X1  _2608_
timestamp 1596033377
transform 1 0 2184 0 -1 610
box -4 -6 52 206
use INVX1  _2594_
timestamp 1596033377
transform -1 0 2264 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert185
timestamp 1596033377
transform -1 0 2312 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert286
timestamp 1596033377
transform 1 0 2312 0 -1 610
box -4 -6 52 206
use INVX1  _2891_
timestamp 1596033377
transform 1 0 2360 0 -1 610
box -4 -6 36 206
use NAND2X1  _2892_
timestamp 1596033377
transform 1 0 2392 0 -1 610
box -4 -6 52 206
use NAND2X1  _2890_
timestamp 1596033377
transform 1 0 2440 0 -1 610
box -4 -6 52 206
use OAI22X1  _2913_
timestamp 1596033377
transform -1 0 2568 0 -1 610
box -4 -6 84 206
use INVX1  _2889_
timestamp 1596033377
transform -1 0 2600 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert156
timestamp 1596033377
transform -1 0 2648 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert85
timestamp 1596033377
transform -1 0 2696 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert183
timestamp 1596033377
transform -1 0 2744 0 -1 610
box -4 -6 52 206
use NAND2X1  _2885_
timestamp 1596033377
transform -1 0 2792 0 -1 610
box -4 -6 52 206
use AOI22X1  _2884_
timestamp 1596033377
transform -1 0 2872 0 -1 610
box -4 -6 84 206
use INVX1  _2882_
timestamp 1596033377
transform 1 0 2872 0 -1 610
box -4 -6 36 206
use INVX1  _2879_
timestamp 1596033377
transform 1 0 2904 0 -1 610
box -4 -6 36 206
use AOI22X1  _2881_
timestamp 1596033377
transform 1 0 3000 0 -1 610
box -4 -6 84 206
use FILL  SFILL29360x4100
timestamp 1596033377
transform -1 0 2952 0 -1 610
box -4 -6 20 206
use FILL  SFILL29520x4100
timestamp 1596033377
transform -1 0 2968 0 -1 610
box -4 -6 20 206
use FILL  SFILL29680x4100
timestamp 1596033377
transform -1 0 2984 0 -1 610
box -4 -6 20 206
use FILL  SFILL29840x4100
timestamp 1596033377
transform -1 0 3000 0 -1 610
box -4 -6 20 206
use INVX1  _2880_
timestamp 1596033377
transform -1 0 3112 0 -1 610
box -4 -6 36 206
use BUFX2  BUFX2_insert84
timestamp 1596033377
transform -1 0 3160 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _4444_
timestamp 1596033377
transform -1 0 3352 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _4445_
timestamp 1596033377
transform -1 0 3544 0 -1 610
box -4 -6 196 206
use AND2X2  _3413_
timestamp 1596033377
transform -1 0 3608 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _3420_
timestamp 1596033377
transform -1 0 3800 0 -1 610
box -4 -6 196 206
use INVX1  _3415_
timestamp 1596033377
transform -1 0 3832 0 -1 610
box -4 -6 36 206
use INVX1  _3407_
timestamp 1596033377
transform 1 0 3832 0 -1 610
box -4 -6 36 206
use NOR2X1  _3412_
timestamp 1596033377
transform -1 0 3912 0 -1 610
box -4 -6 52 206
use OAI21X1  _3387_
timestamp 1596033377
transform -1 0 3976 0 -1 610
box -4 -6 68 206
use NOR2X1  _3416_
timestamp 1596033377
transform 1 0 3976 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _3417_
timestamp 1596033377
transform 1 0 4024 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _3418_
timestamp 1596033377
transform -1 0 4408 0 -1 610
box -4 -6 196 206
use FILL  SFILL44080x4100
timestamp 1596033377
transform -1 0 4424 0 -1 610
box -4 -6 20 206
use BUFX2  _2113_
timestamp 1596033377
transform 1 0 4472 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _3634_
timestamp 1596033377
transform -1 0 4712 0 -1 610
box -4 -6 196 206
use FILL  SFILL44240x4100
timestamp 1596033377
transform -1 0 4440 0 -1 610
box -4 -6 20 206
use FILL  SFILL44400x4100
timestamp 1596033377
transform -1 0 4456 0 -1 610
box -4 -6 20 206
use FILL  SFILL44560x4100
timestamp 1596033377
transform -1 0 4472 0 -1 610
box -4 -6 20 206
use NAND2X1  _3593_
timestamp 1596033377
transform 1 0 4712 0 -1 610
box -4 -6 52 206
use AOI21X1  _3594_
timestamp 1596033377
transform 1 0 4760 0 -1 610
box -4 -6 68 206
use NAND2X1  _3592_
timestamp 1596033377
transform -1 0 4872 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert123
timestamp 1596033377
transform -1 0 4920 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _3633_
timestamp 1596033377
transform -1 0 5112 0 -1 610
box -4 -6 196 206
use NAND2X1  _3620_
timestamp 1596033377
transform 1 0 5112 0 -1 610
box -4 -6 52 206
use AOI21X1  _3621_
timestamp 1596033377
transform 1 0 5160 0 -1 610
box -4 -6 68 206
use BUFX2  BUFX2_insert21
timestamp 1596033377
transform -1 0 5272 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert125
timestamp 1596033377
transform 1 0 5272 0 -1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert20
timestamp 1596033377
transform 1 0 5320 0 -1 610
box -4 -6 52 206
use NAND2X1  _3610_
timestamp 1596033377
transform -1 0 5416 0 -1 610
box -4 -6 52 206
use AOI21X1  _3611_
timestamp 1596033377
transform 1 0 5416 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _3628_
timestamp 1596033377
transform -1 0 5672 0 -1 610
box -4 -6 196 206
use NOR2X1  _3664_
timestamp 1596033377
transform 1 0 5672 0 -1 610
box -4 -6 52 206
use AOI21X1  _3665_
timestamp 1596033377
transform -1 0 5784 0 -1 610
box -4 -6 68 206
use AOI21X1  _3591_
timestamp 1596033377
transform -1 0 5848 0 -1 610
box -4 -6 68 206
use NAND2X1  _3590_
timestamp 1596033377
transform -1 0 5896 0 -1 610
box -4 -6 52 206
use DFFPOSX1  _3640_
timestamp 1596033377
transform 1 0 5960 0 -1 610
box -4 -6 196 206
use FILL  SFILL58960x4100
timestamp 1596033377
transform -1 0 5912 0 -1 610
box -4 -6 20 206
use FILL  SFILL59120x4100
timestamp 1596033377
transform -1 0 5928 0 -1 610
box -4 -6 20 206
use FILL  SFILL59280x4100
timestamp 1596033377
transform -1 0 5944 0 -1 610
box -4 -6 20 206
use FILL  SFILL59440x4100
timestamp 1596033377
transform -1 0 5960 0 -1 610
box -4 -6 20 206
use DFFPOSX1  _4316_
timestamp 1596033377
transform -1 0 6344 0 -1 610
box -4 -6 196 206
use NAND2X1  _3747_
timestamp 1596033377
transform 1 0 6344 0 -1 610
box -4 -6 52 206
use OAI21X1  _3748_
timestamp 1596033377
transform -1 0 6456 0 -1 610
box -4 -6 68 206
use NAND2X1  _3749_
timestamp 1596033377
transform 1 0 6456 0 -1 610
box -4 -6 52 206
use OAI21X1  _3750_
timestamp 1596033377
transform -1 0 6568 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4317_
timestamp 1596033377
transform 1 0 6568 0 -1 610
box -4 -6 196 206
use NAND2X1  _3783_
timestamp 1596033377
transform -1 0 6808 0 -1 610
box -4 -6 52 206
use NAND2X1  _3781_
timestamp 1596033377
transform 1 0 6808 0 -1 610
box -4 -6 52 206
use OAI21X1  _3782_
timestamp 1596033377
transform -1 0 6920 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4348_
timestamp 1596033377
transform -1 0 7112 0 -1 610
box -4 -6 196 206
use OAI21X1  _3776_
timestamp 1596033377
transform 1 0 7112 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _4380_
timestamp 1596033377
transform -1 0 7368 0 -1 610
box -4 -6 196 206
use FILL  FILL71120x4100
timestamp 1596033377
transform -1 0 7384 0 -1 610
box -4 -6 20 206
use FILL  FILL71280x4100
timestamp 1596033377
transform -1 0 7400 0 -1 610
box -4 -6 20 206
use AOI21X1  _2451_
timestamp 1596033377
transform -1 0 72 0 1 610
box -4 -6 68 206
use NAND2X1  _2454_
timestamp 1596033377
transform 1 0 72 0 1 610
box -4 -6 52 206
use NAND3X1  _2535_
timestamp 1596033377
transform -1 0 184 0 1 610
box -4 -6 68 206
use AOI21X1  _2539_
timestamp 1596033377
transform 1 0 184 0 1 610
box -4 -6 68 206
use NOR2X1  _2627_
timestamp 1596033377
transform 1 0 248 0 1 610
box -4 -6 52 206
use OAI21X1  _2629_
timestamp 1596033377
transform 1 0 296 0 1 610
box -4 -6 68 206
use NOR2X1  _2626_
timestamp 1596033377
transform -1 0 408 0 1 610
box -4 -6 52 206
use AOI22X1  _2614_
timestamp 1596033377
transform 1 0 408 0 1 610
box -4 -6 84 206
use NAND2X1  _2615_
timestamp 1596033377
transform 1 0 488 0 1 610
box -4 -6 52 206
use OAI21X1  _2630_
timestamp 1596033377
transform -1 0 600 0 1 610
box -4 -6 68 206
use NOR3X1  _2622_
timestamp 1596033377
transform -1 0 728 0 1 610
box -4 -6 132 206
use BUFX2  BUFX2_insert188
timestamp 1596033377
transform -1 0 776 0 1 610
box -4 -6 52 206
use OR2X2  _2751_
timestamp 1596033377
transform 1 0 776 0 1 610
box -4 -6 68 206
use NAND2X1  _2752_
timestamp 1596033377
transform 1 0 840 0 1 610
box -4 -6 52 206
use AOI22X1  _2755_
timestamp 1596033377
transform 1 0 888 0 1 610
box -4 -6 84 206
use BUFX2  BUFX2_insert301
timestamp 1596033377
transform -1 0 1016 0 1 610
box -4 -6 52 206
use INVX1  _2711_
timestamp 1596033377
transform -1 0 1048 0 1 610
box -4 -6 36 206
use OR2X2  _2753_
timestamp 1596033377
transform -1 0 1112 0 1 610
box -4 -6 68 206
use XNOR2X1  _2933_
timestamp 1596033377
transform -1 0 1224 0 1 610
box -4 -6 116 206
use AND2X2  _2623_
timestamp 1596033377
transform 1 0 1224 0 1 610
box -4 -6 68 206
use NAND2X1  _2538_
timestamp 1596033377
transform -1 0 1336 0 1 610
box -4 -6 52 206
use AOI21X1  _2635_
timestamp 1596033377
transform 1 0 1336 0 1 610
box -4 -6 68 206
use FILL  SFILL14000x6100
timestamp 1596033377
transform 1 0 1400 0 1 610
box -4 -6 20 206
use NAND2X1  _2486_
timestamp 1596033377
transform 1 0 1464 0 1 610
box -4 -6 52 206
use NOR2X1  _2480_
timestamp 1596033377
transform -1 0 1560 0 1 610
box -4 -6 52 206
use NOR2X1  _2537_
timestamp 1596033377
transform 1 0 1560 0 1 610
box -4 -6 52 206
use NOR2X1  _2481_
timestamp 1596033377
transform -1 0 1656 0 1 610
box -4 -6 52 206
use FILL  SFILL14160x6100
timestamp 1596033377
transform 1 0 1416 0 1 610
box -4 -6 20 206
use FILL  SFILL14320x6100
timestamp 1596033377
transform 1 0 1432 0 1 610
box -4 -6 20 206
use FILL  SFILL14480x6100
timestamp 1596033377
transform 1 0 1448 0 1 610
box -4 -6 20 206
use NOR2X1  _2478_
timestamp 1596033377
transform 1 0 1656 0 1 610
box -4 -6 52 206
use INVX1  _2477_
timestamp 1596033377
transform -1 0 1736 0 1 610
box -4 -6 36 206
use XOR2X1  _2536_
timestamp 1596033377
transform -1 0 1848 0 1 610
box -4 -6 116 206
use XNOR2X1  _2483_
timestamp 1596033377
transform 1 0 1848 0 1 610
box -4 -6 116 206
use INVX1  _2809_
timestamp 1596033377
transform -1 0 1992 0 1 610
box -4 -6 36 206
use XNOR2X1  _2482_
timestamp 1596033377
transform -1 0 2104 0 1 610
box -4 -6 116 206
use BUFX2  BUFX2_insert148
timestamp 1596033377
transform -1 0 2152 0 1 610
box -4 -6 52 206
use NAND2X1  _2600_
timestamp 1596033377
transform 1 0 2152 0 1 610
box -4 -6 52 206
use AOI22X1  _2599_
timestamp 1596033377
transform 1 0 2200 0 1 610
box -4 -6 84 206
use BUFX2  BUFX2_insert155
timestamp 1596033377
transform 1 0 2280 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert265
timestamp 1596033377
transform -1 0 2376 0 1 610
box -4 -6 52 206
use INVX1  _2598_
timestamp 1596033377
transform 1 0 2376 0 1 610
box -4 -6 36 206
use NOR2X1  _2894_
timestamp 1596033377
transform -1 0 2456 0 1 610
box -4 -6 52 206
use NAND3X1  _2893_
timestamp 1596033377
transform 1 0 2456 0 1 610
box -4 -6 68 206
use INVX1  _2887_
timestamp 1596033377
transform 1 0 2520 0 1 610
box -4 -6 36 206
use AOI22X1  _2888_
timestamp 1596033377
transform -1 0 2632 0 1 610
box -4 -6 84 206
use INVX1  _2886_
timestamp 1596033377
transform 1 0 2632 0 1 610
box -4 -6 36 206
use OAI21X1  _2914_
timestamp 1596033377
transform 1 0 2664 0 1 610
box -4 -6 68 206
use OAI21X1  _2919_
timestamp 1596033377
transform 1 0 2728 0 1 610
box -4 -6 68 206
use NOR2X1  _2916_
timestamp 1596033377
transform 1 0 2792 0 1 610
box -4 -6 52 206
use INVX1  _2883_
timestamp 1596033377
transform -1 0 2872 0 1 610
box -4 -6 36 206
use AOI21X1  _2918_
timestamp 1596033377
transform 1 0 2872 0 1 610
box -4 -6 68 206
use NAND2X1  _2917_
timestamp 1596033377
transform -1 0 3048 0 1 610
box -4 -6 52 206
use FILL  SFILL29360x6100
timestamp 1596033377
transform 1 0 2936 0 1 610
box -4 -6 20 206
use FILL  SFILL29520x6100
timestamp 1596033377
transform 1 0 2952 0 1 610
box -4 -6 20 206
use FILL  SFILL29680x6100
timestamp 1596033377
transform 1 0 2968 0 1 610
box -4 -6 20 206
use FILL  SFILL29840x6100
timestamp 1596033377
transform 1 0 2984 0 1 610
box -4 -6 20 206
use NOR2X1  _2915_
timestamp 1596033377
transform -1 0 3096 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert147
timestamp 1596033377
transform 1 0 3096 0 1 610
box -4 -6 52 206
use BUFX2  BUFX2_insert158
timestamp 1596033377
transform -1 0 3192 0 1 610
box -4 -6 52 206
use DFFPOSX1  _4431_
timestamp 1596033377
transform -1 0 3384 0 1 610
box -4 -6 196 206
use OAI21X1  _3962_
timestamp 1596033377
transform 1 0 3384 0 1 610
box -4 -6 68 206
use AOI21X1  _3963_
timestamp 1596033377
transform -1 0 3512 0 1 610
box -4 -6 68 206
use DFFPOSX1  _4429_
timestamp 1596033377
transform -1 0 3704 0 1 610
box -4 -6 196 206
use OAI21X1  _3973_
timestamp 1596033377
transform 1 0 3704 0 1 610
box -4 -6 68 206
use AOI21X1  _3974_
timestamp 1596033377
transform -1 0 3832 0 1 610
box -4 -6 68 206
use INVX1  _3528_
timestamp 1596033377
transform 1 0 3832 0 1 610
box -4 -6 36 206
use OAI21X1  _3414_
timestamp 1596033377
transform -1 0 3928 0 1 610
box -4 -6 68 206
use AOI21X1  _3405_
timestamp 1596033377
transform 1 0 3928 0 1 610
box -4 -6 68 206
use OAI21X1  _3403_
timestamp 1596033377
transform 1 0 3992 0 1 610
box -4 -6 68 206
use INVX1  _3535_
timestamp 1596033377
transform -1 0 4088 0 1 610
box -4 -6 36 206
use INVX1  _3402_
timestamp 1596033377
transform -1 0 4120 0 1 610
box -4 -6 36 206
use OAI21X1  _3406_
timestamp 1596033377
transform -1 0 4184 0 1 610
box -4 -6 68 206
use NOR2X1  _3385_
timestamp 1596033377
transform 1 0 4184 0 1 610
box -4 -6 52 206
use OAI21X1  _3386_
timestamp 1596033377
transform 1 0 4232 0 1 610
box -4 -6 68 206
use INVX1  _3388_
timestamp 1596033377
transform 1 0 4296 0 1 610
box -4 -6 36 206
use INVX1  _3521_
timestamp 1596033377
transform 1 0 4328 0 1 610
box -4 -6 36 206
use INVX8  _3563_
timestamp 1596033377
transform 1 0 4360 0 1 610
box -4 -6 84 206
use DFFPOSX1  _3629_
timestamp 1596033377
transform -1 0 4696 0 1 610
box -4 -6 196 206
use FILL  SFILL44400x6100
timestamp 1596033377
transform 1 0 4440 0 1 610
box -4 -6 20 206
use FILL  SFILL44560x6100
timestamp 1596033377
transform 1 0 4456 0 1 610
box -4 -6 20 206
use FILL  SFILL44720x6100
timestamp 1596033377
transform 1 0 4472 0 1 610
box -4 -6 20 206
use FILL  SFILL44880x6100
timestamp 1596033377
transform 1 0 4488 0 1 610
box -4 -6 20 206
use NAND2X1  _3612_
timestamp 1596033377
transform 1 0 4696 0 1 610
box -4 -6 52 206
use AOI21X1  _3613_
timestamp 1596033377
transform -1 0 4808 0 1 610
box -4 -6 68 206
use NAND2X1  _3569_
timestamp 1596033377
transform 1 0 4808 0 1 610
box -4 -6 52 206
use INVX1  _3444_
timestamp 1596033377
transform -1 0 4888 0 1 610
box -4 -6 36 206
use DFFPOSX1  _3632_
timestamp 1596033377
transform -1 0 5080 0 1 610
box -4 -6 196 206
use NAND2X1  _3618_
timestamp 1596033377
transform 1 0 5080 0 1 610
box -4 -6 52 206
use AOI21X1  _3619_
timestamp 1596033377
transform 1 0 5128 0 1 610
box -4 -6 68 206
use INVX1  _3507_
timestamp 1596033377
transform -1 0 5224 0 1 610
box -4 -6 36 206
use AOI21X1  _3579_
timestamp 1596033377
transform -1 0 5288 0 1 610
box -4 -6 68 206
use NAND2X1  _3577_
timestamp 1596033377
transform -1 0 5336 0 1 610
box -4 -6 52 206
use DFFPOSX1  _3642_
timestamp 1596033377
transform 1 0 5336 0 1 610
box -4 -6 196 206
use BUFX2  BUFX2_insert119
timestamp 1596033377
transform -1 0 5576 0 1 610
box -4 -6 52 206
use DFFPOSX1  _4396_
timestamp 1596033377
transform -1 0 5768 0 1 610
box -4 -6 196 206
use AOI21X1  _3884_
timestamp 1596033377
transform 1 0 5768 0 1 610
box -4 -6 68 206
use NOR2X1  _3883_
timestamp 1596033377
transform -1 0 5880 0 1 610
box -4 -6 52 206
use DFFPOSX1  _4333_
timestamp 1596033377
transform 1 0 5944 0 1 610
box -4 -6 196 206
use FILL  SFILL58800x6100
timestamp 1596033377
transform 1 0 5880 0 1 610
box -4 -6 20 206
use FILL  SFILL58960x6100
timestamp 1596033377
transform 1 0 5896 0 1 610
box -4 -6 20 206
use FILL  SFILL59120x6100
timestamp 1596033377
transform 1 0 5912 0 1 610
box -4 -6 20 206
use FILL  SFILL59280x6100
timestamp 1596033377
transform 1 0 5928 0 1 610
box -4 -6 20 206
use BUFX2  BUFX2_insert116
timestamp 1596033377
transform 1 0 6136 0 1 610
box -4 -6 52 206
use MUX2X1  _3972_
timestamp 1596033377
transform 1 0 6184 0 1 610
box -4 -6 100 206
use OAI22X1  _4149_
timestamp 1596033377
transform -1 0 6360 0 1 610
box -4 -6 84 206
use NOR2X1  _4147_
timestamp 1596033377
transform 1 0 6360 0 1 610
box -4 -6 52 206
use OAI21X1  _4148_
timestamp 1596033377
transform -1 0 6472 0 1 610
box -4 -6 68 206
use OAI21X1  _3970_
timestamp 1596033377
transform 1 0 6472 0 1 610
box -4 -6 68 206
use NOR2X1  _3969_
timestamp 1596033377
transform 1 0 6536 0 1 610
box -4 -6 52 206
use OAI22X1  _3971_
timestamp 1596033377
transform 1 0 6584 0 1 610
box -4 -6 84 206
use MUX2X1  _3953_
timestamp 1596033377
transform -1 0 6760 0 1 610
box -4 -6 100 206
use MUX2X1  _4131_
timestamp 1596033377
transform -1 0 6856 0 1 610
box -4 -6 100 206
use MUX2X1  _3964_
timestamp 1596033377
transform 1 0 6856 0 1 610
box -4 -6 100 206
use MUX2X1  _4142_
timestamp 1596033377
transform 1 0 6952 0 1 610
box -4 -6 100 206
use AOI21X1  _3815_
timestamp 1596033377
transform 1 0 7048 0 1 610
box -4 -6 68 206
use NOR2X1  _3814_
timestamp 1596033377
transform 1 0 7112 0 1 610
box -4 -6 52 206
use NOR2X1  _3816_
timestamp 1596033377
transform 1 0 7160 0 1 610
box -4 -6 52 206
use OAI21X1  _3780_
timestamp 1596033377
transform 1 0 7208 0 1 610
box -4 -6 68 206
use AOI21X1  _3817_
timestamp 1596033377
transform -1 0 7336 0 1 610
box -4 -6 68 206
use NOR2X1  _4264_
timestamp 1596033377
transform 1 0 7336 0 1 610
box -4 -6 52 206
use FILL  FILL71280x6100
timestamp 1596033377
transform 1 0 7384 0 1 610
box -4 -6 20 206
use BUFX2  _2104_
timestamp 1596033377
transform -1 0 56 0 -1 1010
box -4 -6 52 206
use XNOR2X1  _2453_
timestamp 1596033377
transform 1 0 56 0 -1 1010
box -4 -6 116 206
use XNOR2X1  _2445_
timestamp 1596033377
transform -1 0 280 0 -1 1010
box -4 -6 116 206
use BUFX2  BUFX2_insert94
timestamp 1596033377
transform -1 0 328 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2628_
timestamp 1596033377
transform -1 0 376 0 -1 1010
box -4 -6 52 206
use INVX1  _2612_
timestamp 1596033377
transform -1 0 408 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert72
timestamp 1596033377
transform -1 0 456 0 -1 1010
box -4 -6 52 206
use INVX1  _2613_
timestamp 1596033377
transform -1 0 488 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert73
timestamp 1596033377
transform 1 0 488 0 -1 1010
box -4 -6 52 206
use INVX1  _2707_
timestamp 1596033377
transform 1 0 536 0 -1 1010
box -4 -6 36 206
use INVX1  _2708_
timestamp 1596033377
transform 1 0 568 0 -1 1010
box -4 -6 36 206
use AOI22X1  _2709_
timestamp 1596033377
transform -1 0 680 0 -1 1010
box -4 -6 84 206
use NAND2X1  _2718_
timestamp 1596033377
transform -1 0 728 0 -1 1010
box -4 -6 52 206
use NOR2X1  _2717_
timestamp 1596033377
transform -1 0 776 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2710_
timestamp 1596033377
transform -1 0 824 0 -1 1010
box -4 -6 52 206
use NAND3X1  _2756_
timestamp 1596033377
transform -1 0 888 0 -1 1010
box -4 -6 68 206
use AOI21X1  _2716_
timestamp 1596033377
transform -1 0 952 0 -1 1010
box -4 -6 68 206
use NOR2X1  _2712_
timestamp 1596033377
transform 1 0 952 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2715_
timestamp 1596033377
transform -1 0 1048 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2714_
timestamp 1596033377
transform 1 0 1048 0 -1 1010
box -4 -6 52 206
use INVX1  _2713_
timestamp 1596033377
transform -1 0 1128 0 -1 1010
box -4 -6 36 206
use BUFX2  BUFX2_insert261
timestamp 1596033377
transform -1 0 1176 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert103
timestamp 1596033377
transform -1 0 1224 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert262
timestamp 1596033377
transform -1 0 1272 0 -1 1010
box -4 -6 52 206
use OAI21X1  _2912_
timestamp 1596033377
transform -1 0 1336 0 -1 1010
box -4 -6 68 206
use XNOR2X1  _2476_
timestamp 1596033377
transform 1 0 1336 0 -1 1010
box -4 -6 116 206
use XNOR2X1  _2475_
timestamp 1596033377
transform 1 0 1512 0 -1 1010
box -4 -6 116 206
use FILL  SFILL14480x8100
timestamp 1596033377
transform -1 0 1464 0 -1 1010
box -4 -6 20 206
use FILL  SFILL14640x8100
timestamp 1596033377
transform -1 0 1480 0 -1 1010
box -4 -6 20 206
use FILL  SFILL14800x8100
timestamp 1596033377
transform -1 0 1496 0 -1 1010
box -4 -6 20 206
use FILL  SFILL14960x8100
timestamp 1596033377
transform -1 0 1512 0 -1 1010
box -4 -6 20 206
use XNOR2X1  _2201_
timestamp 1596033377
transform -1 0 1736 0 -1 1010
box -4 -6 116 206
use NOR2X1  _2935_
timestamp 1596033377
transform 1 0 1736 0 -1 1010
box -4 -6 52 206
use NAND2X1  _2934_
timestamp 1596033377
transform -1 0 1832 0 -1 1010
box -4 -6 52 206
use XNOR2X1  _2932_
timestamp 1596033377
transform 1 0 1832 0 -1 1010
box -4 -6 116 206
use BUFX2  BUFX2_insert239
timestamp 1596033377
transform -1 0 1992 0 -1 1010
box -4 -6 52 206
use NOR2X1  _2303_
timestamp 1596033377
transform 1 0 1992 0 -1 1010
box -4 -6 52 206
use AND2X2  _2304_
timestamp 1596033377
transform -1 0 2104 0 -1 1010
box -4 -6 68 206
use INVX1  _2597_
timestamp 1596033377
transform 1 0 2104 0 -1 1010
box -4 -6 36 206
use AND2X2  _2936_
timestamp 1596033377
transform 1 0 2136 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert290
timestamp 1596033377
transform -1 0 2248 0 -1 1010
box -4 -6 52 206
use AOI21X1  _2920_
timestamp 1596033377
transform 1 0 2248 0 -1 1010
box -4 -6 68 206
use NOR3X1  _2757_
timestamp 1596033377
transform -1 0 2440 0 -1 1010
box -4 -6 132 206
use NOR2X1  _2703_
timestamp 1596033377
transform -1 0 2488 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert289
timestamp 1596033377
transform -1 0 2536 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert241
timestamp 1596033377
transform 1 0 2536 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert57
timestamp 1596033377
transform 1 0 2584 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert288
timestamp 1596033377
transform -1 0 2680 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _4428_
timestamp 1596033377
transform -1 0 2872 0 -1 1010
box -4 -6 196 206
use BUFX2  BUFX2_insert240
timestamp 1596033377
transform 1 0 2872 0 -1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert186
timestamp 1596033377
transform -1 0 3032 0 -1 1010
box -4 -6 52 206
use FILL  SFILL29200x8100
timestamp 1596033377
transform -1 0 2936 0 -1 1010
box -4 -6 20 206
use FILL  SFILL29360x8100
timestamp 1596033377
transform -1 0 2952 0 -1 1010
box -4 -6 20 206
use FILL  SFILL29520x8100
timestamp 1596033377
transform -1 0 2968 0 -1 1010
box -4 -6 20 206
use FILL  SFILL29680x8100
timestamp 1596033377
transform -1 0 2984 0 -1 1010
box -4 -6 20 206
use DFFPOSX1  _4447_
timestamp 1596033377
transform -1 0 3224 0 -1 1010
box -4 -6 196 206
use DFFPOSX1  _4424_
timestamp 1596033377
transform -1 0 3416 0 -1 1010
box -4 -6 196 206
use OAI21X1  _4140_
timestamp 1596033377
transform -1 0 3480 0 -1 1010
box -4 -6 68 206
use AOI21X1  _4141_
timestamp 1596033377
transform -1 0 3544 0 -1 1010
box -4 -6 68 206
use BUFX2  _2089_
timestamp 1596033377
transform 1 0 3544 0 -1 1010
box -4 -6 52 206
use OAI21X1  _4151_
timestamp 1596033377
transform 1 0 3592 0 -1 1010
box -4 -6 68 206
use AOI21X1  _4152_
timestamp 1596033377
transform -1 0 3720 0 -1 1010
box -4 -6 68 206
use INVX1  _3392_
timestamp 1596033377
transform 1 0 3720 0 -1 1010
box -4 -6 36 206
use NAND3X1  _3404_
timestamp 1596033377
transform 1 0 3752 0 -1 1010
box -4 -6 68 206
use AOI22X1  _3396_
timestamp 1596033377
transform 1 0 3816 0 -1 1010
box -4 -6 84 206
use NOR2X1  _3383_
timestamp 1596033377
transform -1 0 3944 0 -1 1010
box -4 -6 52 206
use INVX1  _3384_
timestamp 1596033377
transform -1 0 3976 0 -1 1010
box -4 -6 36 206
use OAI21X1  _3398_
timestamp 1596033377
transform -1 0 4040 0 -1 1010
box -4 -6 68 206
use NOR2X1  _3397_
timestamp 1596033377
transform 1 0 4040 0 -1 1010
box -4 -6 52 206
use NOR2X1  _3390_
timestamp 1596033377
transform 1 0 4088 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3391_
timestamp 1596033377
transform -1 0 4184 0 -1 1010
box -4 -6 52 206
use OAI21X1  _3400_
timestamp 1596033377
transform 1 0 4184 0 -1 1010
box -4 -6 68 206
use INVX1  _3408_
timestamp 1596033377
transform 1 0 4248 0 -1 1010
box -4 -6 36 206
use DFFPOSX1  _3631_
timestamp 1596033377
transform -1 0 4472 0 -1 1010
box -4 -6 196 206
use NAND2X1  _3623_
timestamp 1596033377
transform 1 0 4536 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3624_
timestamp 1596033377
transform 1 0 4584 0 -1 1010
box -4 -6 68 206
use FILL  SFILL44720x8100
timestamp 1596033377
transform -1 0 4488 0 -1 1010
box -4 -6 20 206
use FILL  SFILL44880x8100
timestamp 1596033377
transform -1 0 4504 0 -1 1010
box -4 -6 20 206
use FILL  SFILL45040x8100
timestamp 1596033377
transform -1 0 4520 0 -1 1010
box -4 -6 20 206
use FILL  SFILL45200x8100
timestamp 1596033377
transform -1 0 4536 0 -1 1010
box -4 -6 20 206
use AOI21X1  _3617_
timestamp 1596033377
transform -1 0 4712 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3616_
timestamp 1596033377
transform -1 0 4760 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3622_
timestamp 1596033377
transform -1 0 4808 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3575_
timestamp 1596033377
transform 1 0 4808 0 -1 1010
box -4 -6 52 206
use AOI21X1  _3576_
timestamp 1596033377
transform -1 0 4920 0 -1 1010
box -4 -6 68 206
use AOI21X1  _3570_
timestamp 1596033377
transform -1 0 4984 0 -1 1010
box -4 -6 68 206
use NAND2X1  _3568_
timestamp 1596033377
transform -1 0 5032 0 -1 1010
box -4 -6 52 206
use NAND2X1  _3574_
timestamp 1596033377
transform -1 0 5080 0 -1 1010
box -4 -6 52 206
use MUX2X1  _3961_
timestamp 1596033377
transform -1 0 5176 0 -1 1010
box -4 -6 100 206
use OAI22X1  _3960_
timestamp 1596033377
transform 1 0 5176 0 -1 1010
box -4 -6 84 206
use OAI21X1  _3959_
timestamp 1596033377
transform -1 0 5320 0 -1 1010
box -4 -6 68 206
use MUX2X1  _4139_
timestamp 1596033377
transform -1 0 5416 0 -1 1010
box -4 -6 100 206
use NOR2X1  _4136_
timestamp 1596033377
transform 1 0 5416 0 -1 1010
box -4 -6 52 206
use OAI22X1  _4138_
timestamp 1596033377
transform 1 0 5464 0 -1 1010
box -4 -6 84 206
use MUX2X1  _3957_
timestamp 1596033377
transform -1 0 5640 0 -1 1010
box -4 -6 100 206
use MUX2X1  _4135_
timestamp 1596033377
transform -1 0 5736 0 -1 1010
box -4 -6 100 206
use DFFPOSX1  _4303_
timestamp 1596033377
transform -1 0 5928 0 -1 1010
box -4 -6 196 206
use OAI21X1  _3955_
timestamp 1596033377
transform 1 0 5992 0 -1 1010
box -4 -6 68 206
use FILL  SFILL59280x8100
timestamp 1596033377
transform -1 0 5944 0 -1 1010
box -4 -6 20 206
use FILL  SFILL59440x8100
timestamp 1596033377
transform -1 0 5960 0 -1 1010
box -4 -6 20 206
use FILL  SFILL59600x8100
timestamp 1596033377
transform -1 0 5976 0 -1 1010
box -4 -6 20 206
use FILL  SFILL59760x8100
timestamp 1596033377
transform -1 0 5992 0 -1 1010
box -4 -6 20 206
use OAI22X1  _3956_
timestamp 1596033377
transform 1 0 6056 0 -1 1010
box -4 -6 84 206
use NOR2X1  _4132_
timestamp 1596033377
transform 1 0 6136 0 -1 1010
box -4 -6 52 206
use OAI22X1  _4134_
timestamp 1596033377
transform 1 0 6184 0 -1 1010
box -4 -6 84 206
use OAI21X1  _4133_
timestamp 1596033377
transform -1 0 6328 0 -1 1010
box -4 -6 68 206
use MUX2X1  _4150_
timestamp 1596033377
transform -1 0 6424 0 -1 1010
box -4 -6 100 206
use OAI21X1  _4144_
timestamp 1596033377
transform 1 0 6424 0 -1 1010
box -4 -6 68 206
use OAI22X1  _4145_
timestamp 1596033377
transform -1 0 6568 0 -1 1010
box -4 -6 84 206
use NOR2X1  _4143_
timestamp 1596033377
transform -1 0 6616 0 -1 1010
box -4 -6 52 206
use OAI21X1  _3966_
timestamp 1596033377
transform 1 0 6616 0 -1 1010
box -4 -6 68 206
use OAI22X1  _3967_
timestamp 1596033377
transform -1 0 6760 0 -1 1010
box -4 -6 84 206
use NOR2X1  _3965_
timestamp 1596033377
transform 1 0 6760 0 -1 1010
box -4 -6 52 206
use MUX2X1  _3968_
timestamp 1596033377
transform 1 0 6808 0 -1 1010
box -4 -6 100 206
use MUX2X1  _4146_
timestamp 1596033377
transform 1 0 6904 0 -1 1010
box -4 -6 100 206
use NAND2X1  _3785_
timestamp 1596033377
transform -1 0 7048 0 -1 1010
box -4 -6 52 206
use DFFPOSX1  _4413_
timestamp 1596033377
transform -1 0 7240 0 -1 1010
box -4 -6 196 206
use AOI21X1  _4265_
timestamp 1596033377
transform 1 0 7240 0 -1 1010
box -4 -6 68 206
use NOR2X1  _3818_
timestamp 1596033377
transform -1 0 7352 0 -1 1010
box -4 -6 52 206
use FILL  FILL70960x8100
timestamp 1596033377
transform -1 0 7368 0 -1 1010
box -4 -6 20 206
use FILL  FILL71120x8100
timestamp 1596033377
transform -1 0 7384 0 -1 1010
box -4 -6 20 206
use FILL  FILL71280x8100
timestamp 1596033377
transform -1 0 7400 0 -1 1010
box -4 -6 20 206
use BUFX2  _2105_
timestamp 1596033377
transform -1 0 56 0 1 1010
box -4 -6 52 206
use XNOR2X1  _2452_
timestamp 1596033377
transform -1 0 168 0 1 1010
box -4 -6 116 206
use OAI21X1  _2541_
timestamp 1596033377
transform -1 0 232 0 1 1010
box -4 -6 68 206
use NOR2X1  _2175_
timestamp 1596033377
transform 1 0 232 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert249
timestamp 1596033377
transform -1 0 328 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert248
timestamp 1596033377
transform -1 0 376 0 1 1010
box -4 -6 52 206
use INVX1  _2609_
timestamp 1596033377
transform 1 0 376 0 1 1010
box -4 -6 36 206
use AOI22X1  _2611_
timestamp 1596033377
transform 1 0 408 0 1 1010
box -4 -6 84 206
use AOI22X1  _2706_
timestamp 1596033377
transform 1 0 488 0 1 1010
box -4 -6 84 206
use INVX1  _2705_
timestamp 1596033377
transform -1 0 600 0 1 1010
box -4 -6 36 206
use NOR2X1  _2719_
timestamp 1596033377
transform -1 0 648 0 1 1010
box -4 -6 52 206
use INVX1  _2899_
timestamp 1596033377
transform 1 0 648 0 1 1010
box -4 -6 36 206
use AOI21X1  _2720_
timestamp 1596033377
transform 1 0 680 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert189
timestamp 1596033377
transform 1 0 744 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert98
timestamp 1596033377
transform -1 0 840 0 1 1010
box -4 -6 52 206
use OAI21X1  _2721_
timestamp 1596033377
transform -1 0 904 0 1 1010
box -4 -6 68 206
use NAND2X1  _2754_
timestamp 1596033377
transform 1 0 904 0 1 1010
box -4 -6 52 206
use NOR2X1  _2909_
timestamp 1596033377
transform -1 0 1000 0 1 1010
box -4 -6 52 206
use AOI22X1  _2900_
timestamp 1596033377
transform -1 0 1080 0 1 1010
box -4 -6 84 206
use INVX1  _2896_
timestamp 1596033377
transform 1 0 1080 0 1 1010
box -4 -6 36 206
use NAND2X1  _2910_
timestamp 1596033377
transform 1 0 1112 0 1 1010
box -4 -6 52 206
use AOI21X1  _2911_
timestamp 1596033377
transform 1 0 1160 0 1 1010
box -4 -6 68 206
use NOR2X1  _2908_
timestamp 1596033377
transform 1 0 1224 0 1 1010
box -4 -6 52 206
use INVX1  _2895_
timestamp 1596033377
transform 1 0 1272 0 1 1010
box -4 -6 36 206
use NAND2X1  _2901_
timestamp 1596033377
transform -1 0 1352 0 1 1010
box -4 -6 52 206
use AOI22X1  _2897_
timestamp 1596033377
transform -1 0 1432 0 1 1010
box -4 -6 84 206
use INVX1  _2898_
timestamp 1596033377
transform -1 0 1528 0 1 1010
box -4 -6 36 206
use NOR2X1  _2276_
timestamp 1596033377
transform 1 0 1528 0 1 1010
box -4 -6 52 206
use NOR2X1  _2204_
timestamp 1596033377
transform -1 0 1624 0 1 1010
box -4 -6 52 206
use FILL  SFILL14320x10100
timestamp 1596033377
transform 1 0 1432 0 1 1010
box -4 -6 20 206
use FILL  SFILL14480x10100
timestamp 1596033377
transform 1 0 1448 0 1 1010
box -4 -6 20 206
use FILL  SFILL14640x10100
timestamp 1596033377
transform 1 0 1464 0 1 1010
box -4 -6 20 206
use FILL  SFILL14800x10100
timestamp 1596033377
transform 1 0 1480 0 1 1010
box -4 -6 20 206
use XNOR2X1  _2275_
timestamp 1596033377
transform 1 0 1624 0 1 1010
box -4 -6 116 206
use NAND2X1  _2184_
timestamp 1596033377
transform -1 0 1784 0 1 1010
box -4 -6 52 206
use OR2X2  _2183_
timestamp 1596033377
transform -1 0 1848 0 1 1010
box -4 -6 68 206
use NAND2X1  _2182_
timestamp 1596033377
transform -1 0 1896 0 1 1010
box -4 -6 52 206
use NOR2X1  _2187_
timestamp 1596033377
transform 1 0 1896 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert238
timestamp 1596033377
transform -1 0 1992 0 1 1010
box -4 -6 52 206
use NOR2X1  _2305_
timestamp 1596033377
transform 1 0 1992 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert169
timestamp 1596033377
transform 1 0 2040 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert149
timestamp 1596033377
transform -1 0 2136 0 1 1010
box -4 -6 52 206
use AND2X2  _2193_
timestamp 1596033377
transform -1 0 2200 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert300
timestamp 1596033377
transform -1 0 2248 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert266
timestamp 1596033377
transform -1 0 2296 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert150
timestamp 1596033377
transform -1 0 2344 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert187
timestamp 1596033377
transform 1 0 2344 0 1 1010
box -4 -6 52 206
use OR2X2  _2190_
timestamp 1596033377
transform -1 0 2456 0 1 1010
box -4 -6 68 206
use AOI21X1  _2729_
timestamp 1596033377
transform 1 0 2456 0 1 1010
box -4 -6 68 206
use BUFX2  BUFX2_insert184
timestamp 1596033377
transform -1 0 2568 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert250
timestamp 1596033377
transform -1 0 2616 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert264
timestamp 1596033377
transform -1 0 2664 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _4441_
timestamp 1596033377
transform -1 0 2856 0 1 1010
box -4 -6 196 206
use OAI21X1  _3995_
timestamp 1596033377
transform -1 0 2920 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _4446_
timestamp 1596033377
transform -1 0 3176 0 1 1010
box -4 -6 196 206
use FILL  SFILL29200x10100
timestamp 1596033377
transform 1 0 2920 0 1 1010
box -4 -6 20 206
use FILL  SFILL29360x10100
timestamp 1596033377
transform 1 0 2936 0 1 1010
box -4 -6 20 206
use FILL  SFILL29520x10100
timestamp 1596033377
transform 1 0 2952 0 1 1010
box -4 -6 20 206
use FILL  SFILL29680x10100
timestamp 1596033377
transform 1 0 2968 0 1 1010
box -4 -6 20 206
use AOI21X1  _3996_
timestamp 1596033377
transform -1 0 3240 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _4443_
timestamp 1596033377
transform -1 0 3432 0 1 1010
box -4 -6 196 206
use OAI21X1  _4173_
timestamp 1596033377
transform -1 0 3496 0 1 1010
box -4 -6 68 206
use AOI21X1  _4174_
timestamp 1596033377
transform -1 0 3560 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _4430_
timestamp 1596033377
transform -1 0 3752 0 1 1010
box -4 -6 196 206
use BUFX2  BUFX2_insert136
timestamp 1596033377
transform -1 0 3800 0 1 1010
box -4 -6 52 206
use INVX1  _3393_
timestamp 1596033377
transform 1 0 3800 0 1 1010
box -4 -6 36 206
use NOR2X1  _3394_
timestamp 1596033377
transform -1 0 3880 0 1 1010
box -4 -6 52 206
use NAND2X1  _3395_
timestamp 1596033377
transform -1 0 3928 0 1 1010
box -4 -6 52 206
use AOI21X1  _3409_
timestamp 1596033377
transform 1 0 3928 0 1 1010
box -4 -6 68 206
use INVX1  _3411_
timestamp 1596033377
transform 1 0 3992 0 1 1010
box -4 -6 36 206
use NAND2X1  _3389_
timestamp 1596033377
transform -1 0 4072 0 1 1010
box -4 -6 52 206
use NAND3X1  _3401_
timestamp 1596033377
transform -1 0 4136 0 1 1010
box -4 -6 68 206
use NAND2X1  _3399_
timestamp 1596033377
transform 1 0 4136 0 1 1010
box -4 -6 52 206
use NOR2X1  _3410_
timestamp 1596033377
transform 1 0 4184 0 1 1010
box -4 -6 52 206
use NAND3X1  _3487_
timestamp 1596033377
transform -1 0 4296 0 1 1010
box -4 -6 68 206
use NAND3X1  _3459_
timestamp 1596033377
transform -1 0 4360 0 1 1010
box -4 -6 68 206
use NAND3X1  _3522_
timestamp 1596033377
transform 1 0 4360 0 1 1010
box -4 -6 68 206
use INVX1  _3486_
timestamp 1596033377
transform -1 0 4520 0 1 1010
box -4 -6 36 206
use INVX1  _3451_
timestamp 1596033377
transform 1 0 4520 0 1 1010
box -4 -6 36 206
use NAND3X1  _3480_
timestamp 1596033377
transform -1 0 4616 0 1 1010
box -4 -6 68 206
use NAND3X1  _3515_
timestamp 1596033377
transform -1 0 4680 0 1 1010
box -4 -6 68 206
use FILL  SFILL44240x10100
timestamp 1596033377
transform 1 0 4424 0 1 1010
box -4 -6 20 206
use FILL  SFILL44400x10100
timestamp 1596033377
transform 1 0 4440 0 1 1010
box -4 -6 20 206
use FILL  SFILL44560x10100
timestamp 1596033377
transform 1 0 4456 0 1 1010
box -4 -6 20 206
use FILL  SFILL44720x10100
timestamp 1596033377
transform 1 0 4472 0 1 1010
box -4 -6 20 206
use INVX1  _3465_
timestamp 1596033377
transform -1 0 4712 0 1 1010
box -4 -6 36 206
use NAND3X1  _3473_
timestamp 1596033377
transform -1 0 4776 0 1 1010
box -4 -6 68 206
use INVX1  _3514_
timestamp 1596033377
transform 1 0 4776 0 1 1010
box -4 -6 36 206
use NAND3X1  _3431_
timestamp 1596033377
transform -1 0 4872 0 1 1010
box -4 -6 68 206
use INVX1  _3479_
timestamp 1596033377
transform -1 0 4904 0 1 1010
box -4 -6 36 206
use DFFPOSX1  _3645_
timestamp 1596033377
transform 1 0 4904 0 1 1010
box -4 -6 196 206
use NOR2X1  _3958_
timestamp 1596033377
transform 1 0 5096 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _4335_
timestamp 1596033377
transform 1 0 5144 0 1 1010
box -4 -6 196 206
use AOI21X1  _3888_
timestamp 1596033377
transform 1 0 5336 0 1 1010
box -4 -6 68 206
use NOR2X1  _3887_
timestamp 1596033377
transform -1 0 5448 0 1 1010
box -4 -6 52 206
use OAI21X1  _4137_
timestamp 1596033377
transform 1 0 5448 0 1 1010
box -4 -6 68 206
use OAI21X1  _4170_
timestamp 1596033377
transform 1 0 5512 0 1 1010
box -4 -6 68 206
use OAI22X1  _4171_
timestamp 1596033377
transform -1 0 5656 0 1 1010
box -4 -6 84 206
use OAI21X1  _3992_
timestamp 1596033377
transform 1 0 5656 0 1 1010
box -4 -6 68 206
use NOR2X1  _4169_
timestamp 1596033377
transform -1 0 5768 0 1 1010
box -4 -6 52 206
use OAI22X1  _3993_
timestamp 1596033377
transform -1 0 5848 0 1 1010
box -4 -6 84 206
use NOR2X1  _3991_
timestamp 1596033377
transform 1 0 5848 0 1 1010
box -4 -6 52 206
use MUX2X1  _3994_
timestamp 1596033377
transform -1 0 6056 0 1 1010
box -4 -6 100 206
use FILL  SFILL58960x10100
timestamp 1596033377
transform 1 0 5896 0 1 1010
box -4 -6 20 206
use FILL  SFILL59120x10100
timestamp 1596033377
transform 1 0 5912 0 1 1010
box -4 -6 20 206
use FILL  SFILL59280x10100
timestamp 1596033377
transform 1 0 5928 0 1 1010
box -4 -6 20 206
use FILL  SFILL59440x10100
timestamp 1596033377
transform 1 0 5944 0 1 1010
box -4 -6 20 206
use NAND2X1  _3854_
timestamp 1596033377
transform 1 0 6056 0 1 1010
box -4 -6 52 206
use OAI21X1  _3855_
timestamp 1596033377
transform -1 0 6168 0 1 1010
box -4 -6 68 206
use NOR2X1  _3954_
timestamp 1596033377
transform -1 0 6216 0 1 1010
box -4 -6 52 206
use BUFX2  BUFX2_insert279
timestamp 1596033377
transform 1 0 6216 0 1 1010
box -4 -6 52 206
use DFFPOSX1  _4364_
timestamp 1596033377
transform -1 0 6456 0 1 1010
box -4 -6 196 206
use NAND2X1  _3753_
timestamp 1596033377
transform 1 0 6456 0 1 1010
box -4 -6 52 206
use OAI21X1  _3754_
timestamp 1596033377
transform -1 0 6568 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _4319_
timestamp 1596033377
transform -1 0 6760 0 1 1010
box -4 -6 196 206
use DFFPOSX1  _4365_
timestamp 1596033377
transform -1 0 6952 0 1 1010
box -4 -6 196 206
use OAI21X1  _3786_
timestamp 1596033377
transform 1 0 6952 0 1 1010
box -4 -6 68 206
use DFFPOSX1  _4350_
timestamp 1596033377
transform -1 0 7208 0 1 1010
box -4 -6 196 206
use NOR2X1  _4274_
timestamp 1596033377
transform 1 0 7208 0 1 1010
box -4 -6 52 206
use AOI21X1  _4275_
timestamp 1596033377
transform -1 0 7320 0 1 1010
box -4 -6 68 206
use AOI21X1  _3819_
timestamp 1596033377
transform -1 0 7384 0 1 1010
box -4 -6 68 206
use FILL  FILL71280x10100
timestamp 1596033377
transform 1 0 7384 0 1 1010
box -4 -6 20 206
use OR2X2  _2342_
timestamp 1596033377
transform -1 0 72 0 -1 1410
box -4 -6 68 206
use AND2X2  _2174_
timestamp 1596033377
transform 1 0 72 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert95
timestamp 1596033377
transform -1 0 184 0 -1 1410
box -4 -6 52 206
use INVX1  _2704_
timestamp 1596033377
transform -1 0 216 0 -1 1410
box -4 -6 36 206
use NOR2X1  _2176_
timestamp 1596033377
transform -1 0 264 0 -1 1410
box -4 -6 52 206
use INVX1  _2179_
timestamp 1596033377
transform 1 0 264 0 -1 1410
box -4 -6 36 206
use AOI21X1  _2180_
timestamp 1596033377
transform -1 0 360 0 -1 1410
box -4 -6 68 206
use XNOR2X1  _2177_
timestamp 1596033377
transform -1 0 472 0 -1 1410
box -4 -6 116 206
use INVX1  _2610_
timestamp 1596033377
transform -1 0 504 0 -1 1410
box -4 -6 36 206
use AOI21X1  _2173_
timestamp 1596033377
transform -1 0 568 0 -1 1410
box -4 -6 68 206
use NAND3X1  _2178_
timestamp 1596033377
transform -1 0 632 0 -1 1410
box -4 -6 68 206
use NAND2X1  _2181_
timestamp 1596033377
transform 1 0 632 0 -1 1410
box -4 -6 52 206
use AOI21X1  _2278_
timestamp 1596033377
transform 1 0 680 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert170
timestamp 1596033377
transform -1 0 792 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert104
timestamp 1596033377
transform 1 0 792 0 -1 1410
box -4 -6 52 206
use NAND2X1  _2162_
timestamp 1596033377
transform 1 0 840 0 -1 1410
box -4 -6 52 206
use AND2X2  _2292_
timestamp 1596033377
transform 1 0 888 0 -1 1410
box -4 -6 68 206
use XNOR2X1  _2202_
timestamp 1596033377
transform 1 0 952 0 -1 1410
box -4 -6 116 206
use AOI21X1  _2215_
timestamp 1596033377
transform -1 0 1128 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert263
timestamp 1596033377
transform -1 0 1176 0 -1 1410
box -4 -6 52 206
use INVX1  _2186_
timestamp 1596033377
transform 1 0 1176 0 -1 1410
box -4 -6 36 206
use NAND2X1  _2277_
timestamp 1596033377
transform -1 0 1256 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2274_
timestamp 1596033377
transform 1 0 1256 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2212_
timestamp 1596033377
transform -1 0 1352 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2200_
timestamp 1596033377
transform 1 0 1352 0 -1 1410
box -4 -6 68 206
use AOI21X1  _2206_
timestamp 1596033377
transform 1 0 1480 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2205_
timestamp 1596033377
transform -1 0 1592 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2214_
timestamp 1596033377
transform 1 0 1592 0 -1 1410
box -4 -6 68 206
use FILL  SFILL14160x12100
timestamp 1596033377
transform -1 0 1432 0 -1 1410
box -4 -6 20 206
use FILL  SFILL14320x12100
timestamp 1596033377
transform -1 0 1448 0 -1 1410
box -4 -6 20 206
use FILL  SFILL14480x12100
timestamp 1596033377
transform -1 0 1464 0 -1 1410
box -4 -6 20 206
use FILL  SFILL14640x12100
timestamp 1596033377
transform -1 0 1480 0 -1 1410
box -4 -6 20 206
use XNOR2X1  _2192_
timestamp 1596033377
transform -1 0 1768 0 -1 1410
box -4 -6 116 206
use OAI21X1  _2188_
timestamp 1596033377
transform -1 0 1832 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2208_
timestamp 1596033377
transform -1 0 1880 0 -1 1410
box -4 -6 52 206
use NAND2X1  _2199_
timestamp 1596033377
transform -1 0 1928 0 -1 1410
box -4 -6 52 206
use NOR2X1  _2196_
timestamp 1596033377
transform 1 0 1928 0 -1 1410
box -4 -6 52 206
use AOI21X1  _2195_
timestamp 1596033377
transform 1 0 1976 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2198_
timestamp 1596033377
transform 1 0 2040 0 -1 1410
box -4 -6 52 206
use AND2X2  _2194_
timestamp 1596033377
transform -1 0 2152 0 -1 1410
box -4 -6 68 206
use NOR2X1  _2197_
timestamp 1596033377
transform 1 0 2152 0 -1 1410
box -4 -6 52 206
use NAND2X1  _2191_
timestamp 1596033377
transform -1 0 2248 0 -1 1410
box -4 -6 52 206
use NAND2X1  _2189_
timestamp 1596033377
transform -1 0 2296 0 -1 1410
box -4 -6 52 206
use OR2X2  _2343_
timestamp 1596033377
transform -1 0 2360 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert58
timestamp 1596033377
transform -1 0 2408 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert56
timestamp 1596033377
transform -1 0 2456 0 -1 1410
box -4 -6 52 206
use XOR2X1  _2390_
timestamp 1596033377
transform -1 0 2568 0 -1 1410
box -4 -6 116 206
use NAND2X1  _2410_
timestamp 1596033377
transform 1 0 2568 0 -1 1410
box -4 -6 52 206
use OR2X2  _2411_
timestamp 1596033377
transform 1 0 2616 0 -1 1410
box -4 -6 68 206
use AOI22X1  _2414_
timestamp 1596033377
transform 1 0 2680 0 -1 1410
box -4 -6 84 206
use OAI21X1  _3929_
timestamp 1596033377
transform 1 0 2760 0 -1 1410
box -4 -6 68 206
use AOI21X1  _3930_
timestamp 1596033377
transform -1 0 2888 0 -1 1410
box -4 -6 68 206
use OAI21X1  _3984_
timestamp 1596033377
transform 1 0 2888 0 -1 1410
box -4 -6 68 206
use FILL  SFILL29520x12100
timestamp 1596033377
transform -1 0 2968 0 -1 1410
box -4 -6 20 206
use FILL  SFILL29680x12100
timestamp 1596033377
transform -1 0 2984 0 -1 1410
box -4 -6 20 206
use FILL  SFILL29840x12100
timestamp 1596033377
transform -1 0 3000 0 -1 1410
box -4 -6 20 206
use FILL  SFILL30000x12100
timestamp 1596033377
transform -1 0 3016 0 -1 1410
box -4 -6 20 206
use DFFPOSX1  _4440_
timestamp 1596033377
transform -1 0 3208 0 -1 1410
box -4 -6 196 206
use OAI21X1  _3951_
timestamp 1596033377
transform 1 0 3208 0 -1 1410
box -4 -6 68 206
use AOI21X1  _3952_
timestamp 1596033377
transform -1 0 3336 0 -1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert135
timestamp 1596033377
transform -1 0 3384 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert200
timestamp 1596033377
transform 1 0 3384 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert294
timestamp 1596033377
transform -1 0 3480 0 -1 1410
box -4 -6 52 206
use BUFX2  _2080_
timestamp 1596033377
transform -1 0 3528 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert295
timestamp 1596033377
transform 1 0 3528 0 -1 1410
box -4 -6 52 206
use OAI21X1  _2116_
timestamp 1596033377
transform 1 0 3576 0 -1 1410
box -4 -6 68 206
use BUFX2  _2081_
timestamp 1596033377
transform -1 0 3688 0 -1 1410
box -4 -6 52 206
use INVX1  _3382_
timestamp 1596033377
transform -1 0 3720 0 -1 1410
box -4 -6 36 206
use INVX1  _3916_
timestamp 1596033377
transform -1 0 3752 0 -1 1410
box -4 -6 36 206
use NOR2X1  _3917_
timestamp 1596033377
transform -1 0 3800 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3649_
timestamp 1596033377
transform -1 0 3864 0 -1 1410
box -4 -6 68 206
use AND2X2  _3430_
timestamp 1596033377
transform 1 0 3864 0 -1 1410
box -4 -6 68 206
use NAND3X1  _3529_
timestamp 1596033377
transform 1 0 3928 0 -1 1410
box -4 -6 68 206
use NOR2X1  _3429_
timestamp 1596033377
transform -1 0 4040 0 -1 1410
box -4 -6 52 206
use NAND3X1  _3466_
timestamp 1596033377
transform -1 0 4104 0 -1 1410
box -4 -6 68 206
use INVX1  _3547_
timestamp 1596033377
transform 1 0 4104 0 -1 1410
box -4 -6 36 206
use NOR2X1  _3548_
timestamp 1596033377
transform -1 0 4184 0 -1 1410
box -4 -6 52 206
use INVX4  _3666_
timestamp 1596033377
transform 1 0 4184 0 -1 1410
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert29
timestamp 1596033377
transform -1 0 4376 0 -1 1410
box -4 -6 148 206
use FILL  SFILL43760x12100
timestamp 1596033377
transform -1 0 4392 0 -1 1410
box -4 -6 20 206
use FILL  SFILL43920x12100
timestamp 1596033377
transform -1 0 4408 0 -1 1410
box -4 -6 20 206
use FILL  SFILL44080x12100
timestamp 1596033377
transform -1 0 4424 0 -1 1410
box -4 -6 20 206
use DFFPOSX1  _3625_
timestamp 1596033377
transform -1 0 4632 0 -1 1410
box -4 -6 196 206
use FILL  SFILL44240x12100
timestamp 1596033377
transform -1 0 4440 0 -1 1410
box -4 -6 20 206
use DFFPOSX1  _3641_
timestamp 1596033377
transform 1 0 4632 0 -1 1410
box -4 -6 196 206
use NAND2X1  _3848_
timestamp 1596033377
transform 1 0 4824 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3849_
timestamp 1596033377
transform -1 0 4936 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _4300_
timestamp 1596033377
transform 1 0 4936 0 -1 1410
box -4 -6 196 206
use BUFX2  BUFX2_insert284
timestamp 1596033377
transform -1 0 5176 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert208
timestamp 1596033377
transform -1 0 5224 0 -1 1410
box -4 -6 52 206
use DFFPOSX1  _4412_
timestamp 1596033377
transform 1 0 5224 0 -1 1410
box -4 -6 196 206
use MUX2X1  _3990_
timestamp 1596033377
transform 1 0 5416 0 -1 1410
box -4 -6 100 206
use MUX2X1  _4168_
timestamp 1596033377
transform 1 0 5512 0 -1 1410
box -4 -6 100 206
use MUX2X1  _4172_
timestamp 1596033377
transform -1 0 5704 0 -1 1410
box -4 -6 100 206
use DFFPOSX1  _4399_
timestamp 1596033377
transform -1 0 5896 0 -1 1410
box -4 -6 196 206
use OAI21X1  _3715_
timestamp 1596033377
transform 1 0 5896 0 -1 1410
box -4 -6 68 206
use FILL  SFILL59600x12100
timestamp 1596033377
transform -1 0 5976 0 -1 1410
box -4 -6 20 206
use FILL  SFILL59760x12100
timestamp 1596033377
transform -1 0 5992 0 -1 1410
box -4 -6 20 206
use FILL  SFILL59920x12100
timestamp 1596033377
transform -1 0 6008 0 -1 1410
box -4 -6 20 206
use FILL  SFILL60080x12100
timestamp 1596033377
transform -1 0 6024 0 -1 1410
box -4 -6 20 206
use OAI21X1  _3714_
timestamp 1596033377
transform 1 0 6024 0 -1 1410
box -4 -6 68 206
use OAI22X1  _3989_
timestamp 1596033377
transform -1 0 6168 0 -1 1410
box -4 -6 84 206
use OAI21X1  _3988_
timestamp 1596033377
transform -1 0 6232 0 -1 1410
box -4 -6 68 206
use OAI21X1  _4166_
timestamp 1596033377
transform 1 0 6232 0 -1 1410
box -4 -6 68 206
use OAI22X1  _4167_
timestamp 1596033377
transform 1 0 6296 0 -1 1410
box -4 -6 84 206
use NOR2X1  _4165_
timestamp 1596033377
transform -1 0 6424 0 -1 1410
box -4 -6 52 206
use NOR2X1  _3987_
timestamp 1596033377
transform -1 0 6472 0 -1 1410
box -4 -6 52 206
use OAI21X1  _3716_
timestamp 1596033377
transform 1 0 6472 0 -1 1410
box -4 -6 68 206
use OAI21X1  _3717_
timestamp 1596033377
transform -1 0 6600 0 -1 1410
box -4 -6 68 206
use MUX2X1  _3986_
timestamp 1596033377
transform -1 0 6696 0 -1 1410
box -4 -6 100 206
use MUX2X1  _4164_
timestamp 1596033377
transform -1 0 6792 0 -1 1410
box -4 -6 100 206
use OAI21X1  _3720_
timestamp 1596033377
transform 1 0 6792 0 -1 1410
box -4 -6 68 206
use OAI21X1  _3721_
timestamp 1596033377
transform -1 0 6920 0 -1 1410
box -4 -6 68 206
use DFFPOSX1  _4367_
timestamp 1596033377
transform -1 0 7112 0 -1 1410
box -4 -6 196 206
use DFFPOSX1  _4383_
timestamp 1596033377
transform -1 0 7304 0 -1 1410
box -4 -6 196 206
use NAND2X1  _3779_
timestamp 1596033377
transform -1 0 7352 0 -1 1410
box -4 -6 52 206
use FILL  FILL70960x12100
timestamp 1596033377
transform -1 0 7368 0 -1 1410
box -4 -6 20 206
use FILL  FILL71120x12100
timestamp 1596033377
transform -1 0 7384 0 -1 1410
box -4 -6 20 206
use FILL  FILL71280x12100
timestamp 1596033377
transform -1 0 7400 0 -1 1410
box -4 -6 20 206
use INVX1  _3043_
timestamp 1596033377
transform 1 0 8 0 1 1410
box -4 -6 36 206
use INVX1  _2994_
timestamp 1596033377
transform 1 0 40 0 1 1410
box -4 -6 36 206
use AND2X2  _2358_
timestamp 1596033377
transform 1 0 72 0 1 1410
box -4 -6 68 206
use INVX1  _3046_
timestamp 1596033377
transform 1 0 136 0 1 1410
box -4 -6 36 206
use NOR2X1  _2300_
timestamp 1596033377
transform 1 0 168 0 1 1410
box -4 -6 52 206
use INVX1  _3020_
timestamp 1596033377
transform -1 0 248 0 1 1410
box -4 -6 36 206
use NOR2X1  _2302_
timestamp 1596033377
transform 1 0 248 0 1 1410
box -4 -6 52 206
use AND2X2  _2301_
timestamp 1596033377
transform 1 0 296 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert75
timestamp 1596033377
transform 1 0 360 0 1 1410
box -4 -6 52 206
use NOR2X1  _2170_
timestamp 1596033377
transform -1 0 456 0 1 1410
box -4 -6 52 206
use NOR2X1  _2171_
timestamp 1596033377
transform 1 0 456 0 1 1410
box -4 -6 52 206
use AND2X2  _2169_
timestamp 1596033377
transform -1 0 568 0 1 1410
box -4 -6 68 206
use XOR2X1  _2172_
timestamp 1596033377
transform -1 0 680 0 1 1410
box -4 -6 116 206
use NAND3X1  _3033_
timestamp 1596033377
transform 1 0 680 0 1 1410
box -4 -6 68 206
use NAND3X1  _3059_
timestamp 1596033377
transform 1 0 744 0 1 1410
box -4 -6 68 206
use NAND2X1  _2163_
timestamp 1596033377
transform 1 0 808 0 1 1410
box -4 -6 52 206
use OAI21X1  _2168_
timestamp 1596033377
transform -1 0 920 0 1 1410
box -4 -6 68 206
use NOR2X1  _2165_
timestamp 1596033377
transform -1 0 968 0 1 1410
box -4 -6 52 206
use INVX1  _2164_
timestamp 1596033377
transform 1 0 968 0 1 1410
box -4 -6 36 206
use NOR2X1  _2166_
timestamp 1596033377
transform -1 0 1048 0 1 1410
box -4 -6 52 206
use NAND3X1  _3085_
timestamp 1596033377
transform -1 0 1112 0 1 1410
box -4 -6 68 206
use XNOR2X1  _2185_
timestamp 1596033377
transform 1 0 1112 0 1 1410
box -4 -6 116 206
use INVX1  _3072_
timestamp 1596033377
transform 1 0 1224 0 1 1410
box -4 -6 36 206
use INVX1  _3121_
timestamp 1596033377
transform -1 0 1288 0 1 1410
box -4 -6 36 206
use OR2X2  _2345_
timestamp 1596033377
transform -1 0 1352 0 1 1410
box -4 -6 68 206
use INVX1  _3124_
timestamp 1596033377
transform -1 0 1384 0 1 1410
box -4 -6 36 206
use BUFX2  BUFX2_insert106
timestamp 1596033377
transform 1 0 1384 0 1 1410
box -4 -6 52 206
use AND2X2  _2203_
timestamp 1596033377
transform 1 0 1496 0 1 1410
box -4 -6 68 206
use NAND2X1  _2211_
timestamp 1596033377
transform 1 0 1560 0 1 1410
box -4 -6 52 206
use XNOR2X1  _2210_
timestamp 1596033377
transform 1 0 1608 0 1 1410
box -4 -6 116 206
use FILL  SFILL14320x14100
timestamp 1596033377
transform 1 0 1432 0 1 1410
box -4 -6 20 206
use FILL  SFILL14480x14100
timestamp 1596033377
transform 1 0 1448 0 1 1410
box -4 -6 20 206
use FILL  SFILL14640x14100
timestamp 1596033377
transform 1 0 1464 0 1 1410
box -4 -6 20 206
use FILL  SFILL14800x14100
timestamp 1596033377
transform 1 0 1480 0 1 1410
box -4 -6 20 206
use AOI21X1  _2213_
timestamp 1596033377
transform 1 0 1720 0 1 1410
box -4 -6 68 206
use NOR2X1  _2209_
timestamp 1596033377
transform -1 0 1832 0 1 1410
box -4 -6 52 206
use AND2X2  _2207_
timestamp 1596033377
transform -1 0 1896 0 1 1410
box -4 -6 68 206
use INVX1  _3150_
timestamp 1596033377
transform 1 0 1896 0 1 1410
box -4 -6 36 206
use AND2X2  _2313_
timestamp 1596033377
transform 1 0 1928 0 1 1410
box -4 -6 68 206
use NOR2X1  _2314_
timestamp 1596033377
transform -1 0 2040 0 1 1410
box -4 -6 52 206
use NOR2X1  _2312_
timestamp 1596033377
transform -1 0 2088 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert260
timestamp 1596033377
transform 1 0 2088 0 1 1410
box -4 -6 52 206
use OR2X2  _2344_
timestamp 1596033377
transform 1 0 2136 0 1 1410
box -4 -6 68 206
use INVX1  _3095_
timestamp 1596033377
transform 1 0 2200 0 1 1410
box -4 -6 36 206
use OR2X2  _2346_
timestamp 1596033377
transform 1 0 2232 0 1 1410
box -4 -6 68 206
use INVX1  _3069_
timestamp 1596033377
transform 1 0 2296 0 1 1410
box -4 -6 36 206
use INVX1  _3147_
timestamp 1596033377
transform 1 0 2328 0 1 1410
box -4 -6 36 206
use AND2X2  _2392_
timestamp 1596033377
transform 1 0 2360 0 1 1410
box -4 -6 68 206
use NOR2X1  _2395_
timestamp 1596033377
transform 1 0 2424 0 1 1410
box -4 -6 52 206
use AND2X2  _2394_
timestamp 1596033377
transform 1 0 2472 0 1 1410
box -4 -6 68 206
use OAI22X1  _2396_
timestamp 1596033377
transform -1 0 2616 0 1 1410
box -4 -6 84 206
use BUFX2  BUFX2_insert74
timestamp 1596033377
transform -1 0 2664 0 1 1410
box -4 -6 52 206
use NOR2X1  _2393_
timestamp 1596033377
transform 1 0 2664 0 1 1410
box -4 -6 52 206
use OR2X2  _2413_
timestamp 1596033377
transform -1 0 2776 0 1 1410
box -4 -6 68 206
use NAND2X1  _2412_
timestamp 1596033377
transform 1 0 2776 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert105
timestamp 1596033377
transform -1 0 2872 0 1 1410
box -4 -6 52 206
use DFFPOSX1  _4442_
timestamp 1596033377
transform -1 0 3128 0 1 1410
box -4 -6 196 206
use FILL  SFILL28720x14100
timestamp 1596033377
transform 1 0 2872 0 1 1410
box -4 -6 20 206
use FILL  SFILL28880x14100
timestamp 1596033377
transform 1 0 2888 0 1 1410
box -4 -6 20 206
use FILL  SFILL29040x14100
timestamp 1596033377
transform 1 0 2904 0 1 1410
box -4 -6 20 206
use FILL  SFILL29200x14100
timestamp 1596033377
transform 1 0 2920 0 1 1410
box -4 -6 20 206
use AOI21X1  _3985_
timestamp 1596033377
transform -1 0 3192 0 1 1410
box -4 -6 68 206
use OAI21X1  _3918_
timestamp 1596033377
transform 1 0 3192 0 1 1410
box -4 -6 68 206
use AOI21X1  _3919_
timestamp 1596033377
transform -1 0 3320 0 1 1410
box -4 -6 68 206
use OAI21X1  _4096_
timestamp 1596033377
transform -1 0 3384 0 1 1410
box -4 -6 68 206
use AOI21X1  _4097_
timestamp 1596033377
transform -1 0 3448 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert139
timestamp 1596033377
transform -1 0 3496 0 1 1410
box -4 -6 52 206
use OAI21X1  _2131_
timestamp 1596033377
transform 1 0 3496 0 1 1410
box -4 -6 68 206
use NAND2X1  _2130_
timestamp 1596033377
transform -1 0 3608 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert296
timestamp 1596033377
transform 1 0 3608 0 1 1410
box -4 -6 52 206
use NAND2X1  _2115_
timestamp 1596033377
transform -1 0 3704 0 1 1410
box -4 -6 52 206
use OAI21X1  _2119_
timestamp 1596033377
transform -1 0 3768 0 1 1410
box -4 -6 68 206
use NAND2X1  _2118_
timestamp 1596033377
transform 1 0 3768 0 1 1410
box -4 -6 52 206
use NAND3X1  _3467_
timestamp 1596033377
transform -1 0 3880 0 1 1410
box -4 -6 68 206
use NAND2X1  _3468_
timestamp 1596033377
transform -1 0 3928 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert177
timestamp 1596033377
transform 1 0 3928 0 1 1410
box -4 -6 52 206
use NAND3X1  _3536_
timestamp 1596033377
transform -1 0 4040 0 1 1410
box -4 -6 68 206
use NAND2X1  _3462_
timestamp 1596033377
transform -1 0 4088 0 1 1410
box -4 -6 52 206
use NAND3X1  _3438_
timestamp 1596033377
transform -1 0 4152 0 1 1410
box -4 -6 68 206
use NAND2X1  _3455_
timestamp 1596033377
transform -1 0 4200 0 1 1410
box -4 -6 52 206
use NAND2X1  _3461_
timestamp 1596033377
transform 1 0 4200 0 1 1410
box -4 -6 52 206
use NAND3X1  _3460_
timestamp 1596033377
transform -1 0 4312 0 1 1410
box -4 -6 68 206
use NAND3X1  _3494_
timestamp 1596033377
transform -1 0 4376 0 1 1410
box -4 -6 68 206
use NAND3X1  _3452_
timestamp 1596033377
transform -1 0 4440 0 1 1410
box -4 -6 68 206
use INVX4  _3663_
timestamp 1596033377
transform 1 0 4504 0 1 1410
box -4 -6 52 206
use NAND3X1  _3481_
timestamp 1596033377
transform -1 0 4616 0 1 1410
box -4 -6 68 206
use NAND3X1  _3445_
timestamp 1596033377
transform 1 0 4616 0 1 1410
box -4 -6 68 206
use FILL  SFILL44400x14100
timestamp 1596033377
transform 1 0 4440 0 1 1410
box -4 -6 20 206
use FILL  SFILL44560x14100
timestamp 1596033377
transform 1 0 4456 0 1 1410
box -4 -6 20 206
use FILL  SFILL44720x14100
timestamp 1596033377
transform 1 0 4472 0 1 1410
box -4 -6 20 206
use FILL  SFILL44880x14100
timestamp 1596033377
transform 1 0 4488 0 1 1410
box -4 -6 20 206
use NAND3X1  _3474_
timestamp 1596033377
transform -1 0 4744 0 1 1410
box -4 -6 68 206
use NAND3X1  _3501_
timestamp 1596033377
transform -1 0 4808 0 1 1410
box -4 -6 68 206
use NAND3X1  _3508_
timestamp 1596033377
transform -1 0 4872 0 1 1410
box -4 -6 68 206
use INVX1  _3493_
timestamp 1596033377
transform -1 0 4904 0 1 1410
box -4 -6 36 206
use DFFPOSX1  _4332_
timestamp 1596033377
transform 1 0 4904 0 1 1410
box -4 -6 196 206
use AOI21X1  _3882_
timestamp 1596033377
transform 1 0 5096 0 1 1410
box -4 -6 68 206
use NOR2X1  _3881_
timestamp 1596033377
transform 1 0 5160 0 1 1410
box -4 -6 52 206
use MUX2X1  _4095_
timestamp 1596033377
transform -1 0 5304 0 1 1410
box -4 -6 100 206
use AOI21X1  _4273_
timestamp 1596033377
transform 1 0 5304 0 1 1410
box -4 -6 68 206
use NOR2X1  _4272_
timestamp 1596033377
transform -1 0 5416 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert274
timestamp 1596033377
transform 1 0 5416 0 1 1410
box -4 -6 52 206
use NOR2X1  _4278_
timestamp 1596033377
transform -1 0 5512 0 1 1410
box -4 -6 52 206
use AOI21X1  _4279_
timestamp 1596033377
transform 1 0 5512 0 1 1410
box -4 -6 68 206
use DFFPOSX1  _4415_
timestamp 1596033377
transform -1 0 5768 0 1 1410
box -4 -6 196 206
use NOR2X1  _3673_
timestamp 1596033377
transform 1 0 5768 0 1 1410
box -4 -6 52 206
use AOI21X1  _3674_
timestamp 1596033377
transform -1 0 5880 0 1 1410
box -4 -6 68 206
use BUFX2  BUFX2_insert90
timestamp 1596033377
transform -1 0 5928 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert144
timestamp 1596033377
transform 1 0 5992 0 1 1410
box -4 -6 52 206
use FILL  SFILL59280x14100
timestamp 1596033377
transform 1 0 5928 0 1 1410
box -4 -6 20 206
use FILL  SFILL59440x14100
timestamp 1596033377
transform 1 0 5944 0 1 1410
box -4 -6 20 206
use FILL  SFILL59600x14100
timestamp 1596033377
transform 1 0 5960 0 1 1410
box -4 -6 20 206
use FILL  SFILL59760x14100
timestamp 1596033377
transform 1 0 5976 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_insert93
timestamp 1596033377
transform 1 0 6040 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert211
timestamp 1596033377
transform 1 0 6088 0 1 1410
box -4 -6 52 206
use BUFX2  BUFX2_insert39
timestamp 1596033377
transform 1 0 6136 0 1 1410
box -4 -6 52 206
use OAI22X1  _4090_
timestamp 1596033377
transform -1 0 6264 0 1 1410
box -4 -6 84 206
use NOR2X1  _4088_
timestamp 1596033377
transform -1 0 6312 0 1 1410
box -4 -6 52 206
use OAI21X1  _4089_
timestamp 1596033377
transform 1 0 6312 0 1 1410
box -4 -6 68 206
use MUX2X1  _4086_
timestamp 1596033377
transform -1 0 6472 0 1 1410
box -4 -6 100 206
use MUX2X1  _3906_
timestamp 1596033377
transform 1 0 6472 0 1 1410
box -4 -6 100 206
use MUX2X1  _3975_
timestamp 1596033377
transform -1 0 6664 0 1 1410
box -4 -6 100 206
use MUX2X1  _4153_
timestamp 1596033377
transform -1 0 6760 0 1 1410
box -4 -6 100 206
use DFFPOSX1  _4344_
timestamp 1596033377
transform -1 0 6952 0 1 1410
box -4 -6 196 206
use NAND2X1  _3773_
timestamp 1596033377
transform 1 0 6952 0 1 1410
box -4 -6 52 206
use OAI21X1  _3774_
timestamp 1596033377
transform -1 0 7064 0 1 1410
box -4 -6 68 206
use AOI21X1  _3821_
timestamp 1596033377
transform 1 0 7064 0 1 1410
box -4 -6 68 206
use NOR2X1  _3820_
timestamp 1596033377
transform 1 0 7128 0 1 1410
box -4 -6 52 206
use NOR2X1  _3822_
timestamp 1596033377
transform -1 0 7224 0 1 1410
box -4 -6 52 206
use AOI21X1  _3807_
timestamp 1596033377
transform 1 0 7224 0 1 1410
box -4 -6 68 206
use NOR2X1  _3806_
timestamp 1596033377
transform -1 0 7336 0 1 1410
box -4 -6 52 206
use NAND2X1  _3739_
timestamp 1596033377
transform -1 0 7384 0 1 1410
box -4 -6 52 206
use FILL  FILL71280x14100
timestamp 1596033377
transform 1 0 7384 0 1 1410
box -4 -6 20 206
use INVX1  _2995_
timestamp 1596033377
transform 1 0 8 0 -1 1810
box -4 -6 36 206
use OAI22X1  _2996_
timestamp 1596033377
transform -1 0 120 0 -1 1810
box -4 -6 84 206
use INVX1  _3047_
timestamp 1596033377
transform 1 0 120 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3048_
timestamp 1596033377
transform -1 0 232 0 -1 1810
box -4 -6 84 206
use NOR2X1  _3049_
timestamp 1596033377
transform 1 0 232 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3045_
timestamp 1596033377
transform 1 0 280 0 -1 1810
box -4 -6 84 206
use INVX1  _3044_
timestamp 1596033377
transform -1 0 392 0 -1 1810
box -4 -6 36 206
use INVX1  _2991_
timestamp 1596033377
transform -1 0 424 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3022_
timestamp 1596033377
transform 1 0 424 0 -1 1810
box -4 -6 84 206
use INVX1  _3021_
timestamp 1596033377
transform 1 0 504 0 -1 1810
box -4 -6 36 206
use NOR2X1  _2297_
timestamp 1596033377
transform -1 0 584 0 -1 1810
box -4 -6 52 206
use AND2X2  _2357_
timestamp 1596033377
transform -1 0 648 0 -1 1810
box -4 -6 68 206
use AND2X2  _2298_
timestamp 1596033377
transform 1 0 648 0 -1 1810
box -4 -6 68 206
use AND2X2  _3061_
timestamp 1596033377
transform -1 0 776 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert191
timestamp 1596033377
transform -1 0 824 0 -1 1810
box -4 -6 52 206
use OR2X2  _2340_
timestamp 1596033377
transform -1 0 888 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert299
timestamp 1596033377
transform -1 0 936 0 -1 1810
box -4 -6 52 206
use XNOR2X1  _2167_
timestamp 1596033377
transform -1 0 1048 0 -1 1810
box -4 -6 116 206
use NOR2X1  _3023_
timestamp 1596033377
transform 1 0 1048 0 -1 1810
box -4 -6 52 206
use INVX1  _3018_
timestamp 1596033377
transform 1 0 1096 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3019_
timestamp 1596033377
transform -1 0 1208 0 -1 1810
box -4 -6 84 206
use INVX1  _3017_
timestamp 1596033377
transform -1 0 1240 0 -1 1810
box -4 -6 36 206
use INVX1  _3125_
timestamp 1596033377
transform 1 0 1240 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3126_
timestamp 1596033377
transform -1 0 1352 0 -1 1810
box -4 -6 84 206
use NOR2X1  _3127_
timestamp 1596033377
transform 1 0 1352 0 -1 1810
box -4 -6 52 206
use INVX1  _3122_
timestamp 1596033377
transform 1 0 1400 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3123_
timestamp 1596033377
transform -1 0 1576 0 -1 1810
box -4 -6 84 206
use NOR2X1  _2293_
timestamp 1596033377
transform -1 0 1624 0 -1 1810
box -4 -6 52 206
use FILL  SFILL14320x16100
timestamp 1596033377
transform -1 0 1448 0 -1 1810
box -4 -6 20 206
use FILL  SFILL14480x16100
timestamp 1596033377
transform -1 0 1464 0 -1 1810
box -4 -6 20 206
use FILL  SFILL14640x16100
timestamp 1596033377
transform -1 0 1480 0 -1 1810
box -4 -6 20 206
use FILL  SFILL14800x16100
timestamp 1596033377
transform -1 0 1496 0 -1 1810
box -4 -6 20 206
use NOR2X1  _2291_
timestamp 1596033377
transform 1 0 1624 0 -1 1810
box -4 -6 52 206
use AND2X2  _2310_
timestamp 1596033377
transform 1 0 1672 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2311_
timestamp 1596033377
transform -1 0 1784 0 -1 1810
box -4 -6 52 206
use NOR2X1  _2309_
timestamp 1596033377
transform 1 0 1784 0 -1 1810
box -4 -6 52 206
use AND2X2  _2361_
timestamp 1596033377
transform -1 0 1896 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert81
timestamp 1596033377
transform -1 0 1944 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3074_
timestamp 1596033377
transform 1 0 1944 0 -1 1810
box -4 -6 84 206
use INVX1  _3073_
timestamp 1596033377
transform -1 0 2056 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3152_
timestamp 1596033377
transform 1 0 2056 0 -1 1810
box -4 -6 84 206
use INVX1  _3151_
timestamp 1596033377
transform -1 0 2168 0 -1 1810
box -4 -6 36 206
use OAI22X1  _3100_
timestamp 1596033377
transform 1 0 2168 0 -1 1810
box -4 -6 84 206
use INVX1  _3099_
timestamp 1596033377
transform -1 0 2280 0 -1 1810
box -4 -6 36 206
use OR2X2  _2341_
timestamp 1596033377
transform -1 0 2344 0 -1 1810
box -4 -6 68 206
use OAI22X1  _3071_
timestamp 1596033377
transform 1 0 2344 0 -1 1810
box -4 -6 84 206
use INVX1  _3070_
timestamp 1596033377
transform -1 0 2456 0 -1 1810
box -4 -6 36 206
use NOR2X1  _3075_
timestamp 1596033377
transform -1 0 2504 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3153_
timestamp 1596033377
transform 1 0 2504 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3149_
timestamp 1596033377
transform 1 0 2552 0 -1 1810
box -4 -6 84 206
use INVX1  _3148_
timestamp 1596033377
transform -1 0 2664 0 -1 1810
box -4 -6 36 206
use AND2X2  _2360_
timestamp 1596033377
transform -1 0 2728 0 -1 1810
box -4 -6 68 206
use NOR2X1  _2306_
timestamp 1596033377
transform 1 0 2728 0 -1 1810
box -4 -6 52 206
use AND2X2  _2307_
timestamp 1596033377
transform 1 0 2776 0 -1 1810
box -4 -6 68 206
use XOR2X1  _2372_
timestamp 1596033377
transform 1 0 2840 0 -1 1810
box -4 -6 116 206
use FILL  SFILL29520x16100
timestamp 1596033377
transform -1 0 2968 0 -1 1810
box -4 -6 20 206
use FILL  SFILL29680x16100
timestamp 1596033377
transform -1 0 2984 0 -1 1810
box -4 -6 20 206
use FILL  SFILL29840x16100
timestamp 1596033377
transform -1 0 3000 0 -1 1810
box -4 -6 20 206
use FILL  SFILL30000x16100
timestamp 1596033377
transform -1 0 3016 0 -1 1810
box -4 -6 20 206
use BUFX2  BUFX2_insert298
timestamp 1596033377
transform -1 0 3064 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _4425_
timestamp 1596033377
transform -1 0 3256 0 -1 1810
box -4 -6 196 206
use OAI21X1  _3940_
timestamp 1596033377
transform 1 0 3256 0 -1 1810
box -4 -6 68 206
use AOI21X1  _3941_
timestamp 1596033377
transform -1 0 3384 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert83
timestamp 1596033377
transform -1 0 3432 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert190
timestamp 1596033377
transform -1 0 3480 0 -1 1810
box -4 -6 52 206
use INVX1  _2129_
timestamp 1596033377
transform -1 0 3512 0 -1 1810
box -4 -6 36 206
use DFFPOSX1  _4426_
timestamp 1596033377
transform -1 0 3704 0 -1 1810
box -4 -6 196 206
use OAI21X1  _4118_
timestamp 1596033377
transform -1 0 3768 0 -1 1810
box -4 -6 68 206
use OAI21X1  _4107_
timestamp 1596033377
transform -1 0 3832 0 -1 1810
box -4 -6 68 206
use OAI21X1  _4162_
timestamp 1596033377
transform 1 0 3832 0 -1 1810
box -4 -6 68 206
use AOI21X1  _4163_
timestamp 1596033377
transform -1 0 3960 0 -1 1810
box -4 -6 68 206
use NAND2X1  _4597_
timestamp 1596033377
transform 1 0 3960 0 -1 1810
box -4 -6 52 206
use INVX1  _2114_
timestamp 1596033377
transform -1 0 4040 0 -1 1810
box -4 -6 36 206
use INVX1  _4596_
timestamp 1596033377
transform -1 0 4072 0 -1 1810
box -4 -6 36 206
use NAND2X1  _4585_
timestamp 1596033377
transform 1 0 4072 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3550_
timestamp 1596033377
transform 1 0 4120 0 -1 1810
box -4 -6 52 206
use INVX1  _3549_
timestamp 1596033377
transform -1 0 4200 0 -1 1810
box -4 -6 36 206
use INVX4  _3423_
timestamp 1596033377
transform 1 0 4200 0 -1 1810
box -4 -6 52 206
use INVX1  _3541_
timestamp 1596033377
transform 1 0 4248 0 -1 1810
box -4 -6 36 206
use NOR2X1  _3542_
timestamp 1596033377
transform -1 0 4328 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3434_
timestamp 1596033377
transform -1 0 4376 0 -1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert130
timestamp 1596033377
transform -1 0 4424 0 -1 1810
box -4 -6 52 206
use AND2X2  _3562_
timestamp 1596033377
transform -1 0 4552 0 -1 1810
box -4 -6 68 206
use NOR2X1  _3554_
timestamp 1596033377
transform 1 0 4552 0 -1 1810
box -4 -6 52 206
use INVX1  _3553_
timestamp 1596033377
transform -1 0 4632 0 -1 1810
box -4 -6 36 206
use FILL  SFILL44240x16100
timestamp 1596033377
transform -1 0 4440 0 -1 1810
box -4 -6 20 206
use FILL  SFILL44400x16100
timestamp 1596033377
transform -1 0 4456 0 -1 1810
box -4 -6 20 206
use FILL  SFILL44560x16100
timestamp 1596033377
transform -1 0 4472 0 -1 1810
box -4 -6 20 206
use FILL  SFILL44720x16100
timestamp 1596033377
transform -1 0 4488 0 -1 1810
box -4 -6 20 206
use BUFX2  BUFX2_insert129
timestamp 1596033377
transform 1 0 4632 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3476_
timestamp 1596033377
transform -1 0 4728 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3482_
timestamp 1596033377
transform 1 0 4728 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3469_
timestamp 1596033377
transform 1 0 4776 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3552_
timestamp 1596033377
transform 1 0 4824 0 -1 1810
box -4 -6 52 206
use INVX1  _3551_
timestamp 1596033377
transform -1 0 4904 0 -1 1810
box -4 -6 36 206
use NAND2X1  _3475_
timestamp 1596033377
transform 1 0 4904 0 -1 1810
box -4 -6 52 206
use INVX4  _3672_
timestamp 1596033377
transform -1 0 5000 0 -1 1810
box -4 -6 52 206
use INVX4  _3669_
timestamp 1596033377
transform -1 0 5048 0 -1 1810
box -4 -6 52 206
use DFFPOSX1  _4328_
timestamp 1596033377
transform 1 0 5048 0 -1 1810
box -4 -6 196 206
use OAI21X1  _3913_
timestamp 1596033377
transform 1 0 5240 0 -1 1810
box -4 -6 68 206
use OAI22X1  _3914_
timestamp 1596033377
transform -1 0 5384 0 -1 1810
box -4 -6 84 206
use NOR2X1  _3912_
timestamp 1596033377
transform -1 0 5432 0 -1 1810
box -4 -6 52 206
use MUX2X1  _3915_
timestamp 1596033377
transform -1 0 5528 0 -1 1810
box -4 -6 100 206
use NOR2X1  _4092_
timestamp 1596033377
transform 1 0 5528 0 -1 1810
box -4 -6 52 206
use OAI22X1  _4094_
timestamp 1596033377
transform -1 0 5656 0 -1 1810
box -4 -6 84 206
use OAI21X1  _4093_
timestamp 1596033377
transform 1 0 5656 0 -1 1810
box -4 -6 68 206
use NOR2X1  _3980_
timestamp 1596033377
transform 1 0 5720 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3982_
timestamp 1596033377
transform -1 0 5848 0 -1 1810
box -4 -6 84 206
use OAI21X1  _3981_
timestamp 1596033377
transform 1 0 5848 0 -1 1810
box -4 -6 68 206
use MUX2X1  _3983_
timestamp 1596033377
transform -1 0 6072 0 -1 1810
box -4 -6 100 206
use FILL  SFILL59120x16100
timestamp 1596033377
transform -1 0 5928 0 -1 1810
box -4 -6 20 206
use FILL  SFILL59280x16100
timestamp 1596033377
transform -1 0 5944 0 -1 1810
box -4 -6 20 206
use FILL  SFILL59440x16100
timestamp 1596033377
transform -1 0 5960 0 -1 1810
box -4 -6 20 206
use FILL  SFILL59600x16100
timestamp 1596033377
transform -1 0 5976 0 -1 1810
box -4 -6 20 206
use MUX2X1  _4161_
timestamp 1596033377
transform -1 0 6168 0 -1 1810
box -4 -6 100 206
use BUFX2  BUFX2_insert280
timestamp 1596033377
transform 1 0 6168 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3705_
timestamp 1596033377
transform 1 0 6216 0 -1 1810
box -4 -6 52 206
use NAND2X1  _3738_
timestamp 1596033377
transform -1 0 6312 0 -1 1810
box -4 -6 52 206
use NOR2X1  _3650_
timestamp 1596033377
transform 1 0 6312 0 -1 1810
box -4 -6 52 206
use OAI21X1  _4155_
timestamp 1596033377
transform 1 0 6360 0 -1 1810
box -4 -6 68 206
use OAI22X1  _4156_
timestamp 1596033377
transform -1 0 6504 0 -1 1810
box -4 -6 84 206
use NOR2X1  _4154_
timestamp 1596033377
transform -1 0 6552 0 -1 1810
box -4 -6 52 206
use OAI22X1  _3978_
timestamp 1596033377
transform 1 0 6552 0 -1 1810
box -4 -6 84 206
use NOR2X1  _3976_
timestamp 1596033377
transform 1 0 6632 0 -1 1810
box -4 -6 52 206
use OAI21X1  _3909_
timestamp 1596033377
transform 1 0 6680 0 -1 1810
box -4 -6 68 206
use OAI22X1  _3910_
timestamp 1596033377
transform -1 0 6824 0 -1 1810
box -4 -6 84 206
use NOR2X1  _3908_
timestamp 1596033377
transform -1 0 6872 0 -1 1810
box -4 -6 52 206
use OAI21X1  _3706_
timestamp 1596033377
transform 1 0 6872 0 -1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert6
timestamp 1596033377
transform -1 0 6984 0 -1 1810
box -4 -6 52 206
use AOI21X1  _3835_
timestamp 1596033377
transform 1 0 6984 0 -1 1810
box -4 -6 68 206
use NAND2X1  _3787_
timestamp 1596033377
transform 1 0 7048 0 -1 1810
box -4 -6 52 206
use OAI21X1  _3788_
timestamp 1596033377
transform -1 0 7160 0 -1 1810
box -4 -6 68 206
use DFFPOSX1  _4351_
timestamp 1596033377
transform -1 0 7352 0 -1 1810
box -4 -6 196 206
use FILL  FILL70960x16100
timestamp 1596033377
transform -1 0 7368 0 -1 1810
box -4 -6 20 206
use FILL  FILL71120x16100
timestamp 1596033377
transform -1 0 7384 0 -1 1810
box -4 -6 20 206
use FILL  FILL71280x16100
timestamp 1596033377
transform -1 0 7400 0 -1 1810
box -4 -6 20 206
use NOR2X1  _2997_
timestamp 1596033377
transform -1 0 56 0 1 1810
box -4 -6 52 206
use INVX1  _2992_
timestamp 1596033377
transform 1 0 56 0 1 1810
box -4 -6 36 206
use OAI22X1  _2993_
timestamp 1596033377
transform -1 0 168 0 1 1810
box -4 -6 84 206
use NAND2X1  _3063_
timestamp 1596033377
transform 1 0 168 0 1 1810
box -4 -6 52 206
use NAND3X1  _3068_
timestamp 1596033377
transform -1 0 280 0 1 1810
box -4 -6 68 206
use NOR2X1  _3067_
timestamp 1596033377
transform -1 0 328 0 1 1810
box -4 -6 52 206
use INVX1  _3435_
timestamp 1596033377
transform 1 0 328 0 1 1810
box -4 -6 36 206
use NAND2X1  _3057_
timestamp 1596033377
transform 1 0 360 0 1 1810
box -4 -6 52 206
use NAND3X1  _3062_
timestamp 1596033377
transform 1 0 408 0 1 1810
box -4 -6 68 206
use NAND3X1  _3058_
timestamp 1596033377
transform 1 0 472 0 1 1810
box -4 -6 68 206
use NOR2X1  _2299_
timestamp 1596033377
transform 1 0 536 0 1 1810
box -4 -6 52 206
use AND2X2  _2356_
timestamp 1596033377
transform -1 0 648 0 1 1810
box -4 -6 68 206
use NAND3X1  _3006_
timestamp 1596033377
transform -1 0 712 0 1 1810
box -4 -6 68 206
use NOR2X1  _2294_
timestamp 1596033377
transform -1 0 760 0 1 1810
box -4 -6 52 206
use NOR2X1  _2296_
timestamp 1596033377
transform 1 0 760 0 1 1810
box -4 -6 52 206
use AND2X2  _2295_
timestamp 1596033377
transform -1 0 872 0 1 1810
box -4 -6 68 206
use BUFX2  BUFX2_insert272
timestamp 1596033377
transform 1 0 872 0 1 1810
box -4 -6 52 206
use NAND3X1  _3007_
timestamp 1596033377
transform 1 0 920 0 1 1810
box -4 -6 68 206
use NAND3X1  _3137_
timestamp 1596033377
transform 1 0 984 0 1 1810
box -4 -6 68 206
use AND2X2  _3139_
timestamp 1596033377
transform 1 0 1048 0 1 1810
box -4 -6 68 206
use AND2X2  _3087_
timestamp 1596033377
transform 1 0 1112 0 1 1810
box -4 -6 68 206
use NAND3X1  _3140_
timestamp 1596033377
transform -1 0 1240 0 1 1810
box -4 -6 68 206
use NOR2X1  _3145_
timestamp 1596033377
transform 1 0 1240 0 1 1810
box -4 -6 52 206
use NAND3X1  _3146_
timestamp 1596033377
transform -1 0 1352 0 1 1810
box -4 -6 68 206
use NAND3X1  _3136_
timestamp 1596033377
transform -1 0 1416 0 1 1810
box -4 -6 68 206
use NAND2X1  _3141_
timestamp 1596033377
transform -1 0 1528 0 1 1810
box -4 -6 52 206
use NAND3X1  _2976_
timestamp 1596033377
transform -1 0 1592 0 1 1810
box -4 -6 68 206
use NAND3X1  _3111_
timestamp 1596033377
transform -1 0 1656 0 1 1810
box -4 -6 68 206
use FILL  SFILL14160x18100
timestamp 1596033377
transform 1 0 1416 0 1 1810
box -4 -6 20 206
use FILL  SFILL14320x18100
timestamp 1596033377
transform 1 0 1432 0 1 1810
box -4 -6 20 206
use FILL  SFILL14480x18100
timestamp 1596033377
transform 1 0 1448 0 1 1810
box -4 -6 20 206
use FILL  SFILL14640x18100
timestamp 1596033377
transform 1 0 1464 0 1 1810
box -4 -6 20 206
use NAND3X1  _3163_
timestamp 1596033377
transform -1 0 1720 0 1 1810
box -4 -6 68 206
use AND2X2  _3165_
timestamp 1596033377
transform 1 0 1720 0 1 1810
box -4 -6 68 206
use INVX1  _3449_
timestamp 1596033377
transform 1 0 1784 0 1 1810
box -4 -6 36 206
use NAND3X1  _3162_
timestamp 1596033377
transform -1 0 1880 0 1 1810
box -4 -6 68 206
use NAND3X1  _3084_
timestamp 1596033377
transform -1 0 1944 0 1 1810
box -4 -6 68 206
use NAND3X1  _3088_
timestamp 1596033377
transform -1 0 2008 0 1 1810
box -4 -6 68 206
use NAND2X1  _3083_
timestamp 1596033377
transform -1 0 2056 0 1 1810
box -4 -6 52 206
use NAND3X1  _3166_
timestamp 1596033377
transform -1 0 2120 0 1 1810
box -4 -6 68 206
use NAND2X1  _3161_
timestamp 1596033377
transform -1 0 2168 0 1 1810
box -4 -6 52 206
use NOR2X1  _3093_
timestamp 1596033377
transform 1 0 2168 0 1 1810
box -4 -6 52 206
use NOR2X1  _3101_
timestamp 1596033377
transform 1 0 2216 0 1 1810
box -4 -6 52 206
use OAI22X1  _3097_
timestamp 1596033377
transform 1 0 2264 0 1 1810
box -4 -6 84 206
use INVX1  _3096_
timestamp 1596033377
transform -1 0 2376 0 1 1810
box -4 -6 36 206
use NOR2X1  _3171_
timestamp 1596033377
transform -1 0 2424 0 1 1810
box -4 -6 52 206
use NAND2X1  _3115_
timestamp 1596033377
transform -1 0 2472 0 1 1810
box -4 -6 52 206
use NAND3X1  _3094_
timestamp 1596033377
transform 1 0 2472 0 1 1810
box -4 -6 68 206
use NAND3X1  _3172_
timestamp 1596033377
transform 1 0 2536 0 1 1810
box -4 -6 68 206
use INVX1  _3456_
timestamp 1596033377
transform 1 0 2600 0 1 1810
box -4 -6 36 206
use XNOR2X1  _2418_
timestamp 1596033377
transform 1 0 2632 0 1 1810
box -4 -6 116 206
use NOR2X1  _2308_
timestamp 1596033377
transform 1 0 2744 0 1 1810
box -4 -6 52 206
use INVX1  _3477_
timestamp 1596033377
transform -1 0 2824 0 1 1810
box -4 -6 36 206
use INVX1  _3463_
timestamp 1596033377
transform -1 0 2856 0 1 1810
box -4 -6 36 206
use OAI21X1  _3436_
timestamp 1596033377
transform -1 0 2920 0 1 1810
box -4 -6 68 206
use OAI21X1  _3464_
timestamp 1596033377
transform -1 0 3048 0 1 1810
box -4 -6 68 206
use FILL  SFILL29200x18100
timestamp 1596033377
transform 1 0 2920 0 1 1810
box -4 -6 20 206
use FILL  SFILL29360x18100
timestamp 1596033377
transform 1 0 2936 0 1 1810
box -4 -6 20 206
use FILL  SFILL29520x18100
timestamp 1596033377
transform 1 0 2952 0 1 1810
box -4 -6 20 206
use FILL  SFILL29680x18100
timestamp 1596033377
transform 1 0 2968 0 1 1810
box -4 -6 20 206
use OAI21X1  _3457_
timestamp 1596033377
transform -1 0 3112 0 1 1810
box -4 -6 68 206
use INVX1  _3470_
timestamp 1596033377
transform -1 0 3144 0 1 1810
box -4 -6 36 206
use OAI21X1  _3471_
timestamp 1596033377
transform -1 0 3208 0 1 1810
box -4 -6 68 206
use OAI21X1  _3427_
timestamp 1596033377
transform -1 0 3272 0 1 1810
box -4 -6 68 206
use OAI21X1  _3478_
timestamp 1596033377
transform -1 0 3336 0 1 1810
box -4 -6 68 206
use OAI21X1  _3450_
timestamp 1596033377
transform 1 0 3336 0 1 1810
box -4 -6 68 206
use OAI21X1  _2134_
timestamp 1596033377
transform 1 0 3400 0 1 1810
box -4 -6 68 206
use NAND2X1  _2133_
timestamp 1596033377
transform 1 0 3464 0 1 1810
box -4 -6 52 206
use NAND2X1  _4600_
timestamp 1596033377
transform -1 0 3560 0 1 1810
box -4 -6 52 206
use OAI21X1  _4601_
timestamp 1596033377
transform -1 0 3624 0 1 1810
box -4 -6 68 206
use INVX1  _4599_
timestamp 1596033377
transform -1 0 3656 0 1 1810
box -4 -6 36 206
use NAND2X1  _4603_
timestamp 1596033377
transform -1 0 3704 0 1 1810
box -4 -6 52 206
use AOI21X1  _4119_
timestamp 1596033377
transform -1 0 3768 0 1 1810
box -4 -6 68 206
use AOI21X1  _4108_
timestamp 1596033377
transform -1 0 3832 0 1 1810
box -4 -6 68 206
use NAND2X1  _4582_
timestamp 1596033377
transform 1 0 3832 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert181
timestamp 1596033377
transform -1 0 3928 0 1 1810
box -4 -6 52 206
use OAI21X1  _4598_
timestamp 1596033377
transform -1 0 3992 0 1 1810
box -4 -6 68 206
use OAI21X1  _4583_
timestamp 1596033377
transform -1 0 4056 0 1 1810
box -4 -6 68 206
use INVX1  _4593_
timestamp 1596033377
transform -1 0 4088 0 1 1810
box -4 -6 36 206
use OAI21X1  _4586_
timestamp 1596033377
transform -1 0 4152 0 1 1810
box -4 -6 68 206
use NAND3X1  _3439_
timestamp 1596033377
transform -1 0 4216 0 1 1810
box -4 -6 68 206
use INVX1  _4602_
timestamp 1596033377
transform -1 0 4248 0 1 1810
box -4 -6 36 206
use INVX1  _4584_
timestamp 1596033377
transform -1 0 4280 0 1 1810
box -4 -6 36 206
use NAND2X1  _3440_
timestamp 1596033377
transform -1 0 4328 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_insert176
timestamp 1596033377
transform -1 0 4376 0 1 1810
box -4 -6 52 206
use NAND3X1  _3453_
timestamp 1596033377
transform -1 0 4440 0 1 1810
box -4 -6 68 206
use INVX1  _4581_
timestamp 1596033377
transform -1 0 4536 0 1 1810
box -4 -6 36 206
use NOR2X1  _3540_
timestamp 1596033377
transform 1 0 4536 0 1 1810
box -4 -6 52 206
use INVX1  _3539_
timestamp 1596033377
transform -1 0 4616 0 1 1810
box -4 -6 36 206
use NAND2X1  _3422_
timestamp 1596033377
transform 1 0 4616 0 1 1810
box -4 -6 52 206
use FILL  SFILL44400x18100
timestamp 1596033377
transform 1 0 4440 0 1 1810
box -4 -6 20 206
use FILL  SFILL44560x18100
timestamp 1596033377
transform 1 0 4456 0 1 1810
box -4 -6 20 206
use FILL  SFILL44720x18100
timestamp 1596033377
transform 1 0 4472 0 1 1810
box -4 -6 20 206
use FILL  SFILL44880x18100
timestamp 1596033377
transform 1 0 4488 0 1 1810
box -4 -6 20 206
use NAND2X1  _3433_
timestamp 1596033377
transform 1 0 4664 0 1 1810
box -4 -6 52 206
use NAND3X1  _3432_
timestamp 1596033377
transform -1 0 4776 0 1 1810
box -4 -6 68 206
use NAND3X1  _3509_
timestamp 1596033377
transform 1 0 4776 0 1 1810
box -4 -6 68 206
use INVX4  _3654_
timestamp 1596033377
transform 1 0 4840 0 1 1810
box -4 -6 52 206
use INVX4  _3647_
timestamp 1596033377
transform 1 0 4888 0 1 1810
box -4 -6 52 206
use DFFPOSX1  _4302_
timestamp 1596033377
transform 1 0 4936 0 1 1810
box -4 -6 196 206
use OAI21X1  _3853_
timestamp 1596033377
transform 1 0 5128 0 1 1810
box -4 -6 68 206
use NAND2X1  _3852_
timestamp 1596033377
transform -1 0 5240 0 1 1810
box -4 -6 52 206
use NOR2X1  _3873_
timestamp 1596033377
transform 1 0 5240 0 1 1810
box -4 -6 52 206
use AOI21X1  _3874_
timestamp 1596033377
transform -1 0 5352 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _4398_
timestamp 1596033377
transform 1 0 5352 0 1 1810
box -4 -6 196 206
use NOR2X1  _3670_
timestamp 1596033377
transform 1 0 5544 0 1 1810
box -4 -6 52 206
use AOI21X1  _3671_
timestamp 1596033377
transform -1 0 5656 0 1 1810
box -4 -6 68 206
use OAI21X1  _4159_
timestamp 1596033377
transform 1 0 5656 0 1 1810
box -4 -6 68 206
use NOR2X1  _4158_
timestamp 1596033377
transform 1 0 5720 0 1 1810
box -4 -6 52 206
use MUX2X1  _3979_
timestamp 1596033377
transform 1 0 5768 0 1 1810
box -4 -6 100 206
use OAI22X1  _4160_
timestamp 1596033377
transform 1 0 5864 0 1 1810
box -4 -6 84 206
use MUX2X1  _4157_
timestamp 1596033377
transform 1 0 6008 0 1 1810
box -4 -6 100 206
use FILL  SFILL59440x18100
timestamp 1596033377
transform 1 0 5944 0 1 1810
box -4 -6 20 206
use FILL  SFILL59600x18100
timestamp 1596033377
transform 1 0 5960 0 1 1810
box -4 -6 20 206
use FILL  SFILL59760x18100
timestamp 1596033377
transform 1 0 5976 0 1 1810
box -4 -6 20 206
use FILL  SFILL59920x18100
timestamp 1596033377
transform 1 0 5992 0 1 1810
box -4 -6 20 206
use NOR2X1  _3648_
timestamp 1596033377
transform 1 0 6104 0 1 1810
box -4 -6 52 206
use NOR2X1  _3838_
timestamp 1596033377
transform 1 0 6152 0 1 1810
box -4 -6 52 206
use INVX1  _3699_
timestamp 1596033377
transform 1 0 6200 0 1 1810
box -4 -6 36 206
use NAND2X1  _3704_
timestamp 1596033377
transform -1 0 6280 0 1 1810
box -4 -6 52 206
use NOR2X1  _3701_
timestamp 1596033377
transform 1 0 6280 0 1 1810
box -4 -6 52 206
use INVX1  _3700_
timestamp 1596033377
transform -1 0 6360 0 1 1810
box -4 -6 36 206
use INVX1  _3702_
timestamp 1596033377
transform 1 0 6360 0 1 1810
box -4 -6 36 206
use NOR2X1  _3771_
timestamp 1596033377
transform 1 0 6392 0 1 1810
box -4 -6 52 206
use NAND2X1  _3772_
timestamp 1596033377
transform -1 0 6488 0 1 1810
box -4 -6 52 206
use AND2X2  _3805_
timestamp 1596033377
transform 1 0 6488 0 1 1810
box -4 -6 68 206
use OAI21X1  _3977_
timestamp 1596033377
transform 1 0 6552 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _4414_
timestamp 1596033377
transform -1 0 6808 0 1 1810
box -4 -6 196 206
use NOR2X1  _4276_
timestamp 1596033377
transform 1 0 6808 0 1 1810
box -4 -6 52 206
use AOI21X1  _4277_
timestamp 1596033377
transform -1 0 6920 0 1 1810
box -4 -6 68 206
use OAI21X1  _3707_
timestamp 1596033377
transform -1 0 6984 0 1 1810
box -4 -6 68 206
use DFFPOSX1  _4360_
timestamp 1596033377
transform -1 0 7176 0 1 1810
box -4 -6 196 206
use DFFPOSX1  _4312_
timestamp 1596033377
transform -1 0 7368 0 1 1810
box -4 -6 196 206
use FILL  FILL71120x18100
timestamp 1596033377
transform 1 0 7368 0 1 1810
box -4 -6 20 206
use FILL  FILL71280x18100
timestamp 1596033377
transform 1 0 7384 0 1 1810
box -4 -6 20 206
use NAND3X1  _3016_
timestamp 1596033377
transform 1 0 8 0 -1 2210
box -4 -6 68 206
use AOI22X1  _3065_
timestamp 1596033377
transform -1 0 152 0 -1 2210
box -4 -6 84 206
use NAND3X1  _3066_
timestamp 1596033377
transform -1 0 216 0 -1 2210
box -4 -6 68 206
use NOR2X1  _3056_
timestamp 1596033377
transform -1 0 264 0 -1 2210
box -4 -6 52 206
use NOR2X1  _3015_
timestamp 1596033377
transform 1 0 264 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3011_
timestamp 1596033377
transform -1 0 360 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3031_
timestamp 1596033377
transform 1 0 360 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3036_
timestamp 1596033377
transform 1 0 408 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3032_
timestamp 1596033377
transform -1 0 536 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3037_
timestamp 1596033377
transform -1 0 584 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3005_
timestamp 1596033377
transform 1 0 584 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3010_
timestamp 1596033377
transform 1 0 632 0 -1 2210
box -4 -6 68 206
use AND2X2  _3009_
timestamp 1596033377
transform -1 0 760 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert225
timestamp 1596033377
transform -1 0 808 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert269
timestamp 1596033377
transform 1 0 808 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert66
timestamp 1596033377
transform 1 0 856 0 -1 2210
box -4 -6 52 206
use NAND3X1  _3138_
timestamp 1596033377
transform -1 0 968 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3086_
timestamp 1596033377
transform -1 0 1032 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3112_
timestamp 1596033377
transform -1 0 1096 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3164_
timestamp 1596033377
transform -1 0 1160 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert235
timestamp 1596033377
transform -1 0 1208 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3135_
timestamp 1596033377
transform 1 0 1208 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert214
timestamp 1596033377
transform 1 0 1256 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert228
timestamp 1596033377
transform 1 0 1304 0 -1 2210
box -4 -6 52 206
use AOI22X1  _3143_
timestamp 1596033377
transform 1 0 1352 0 -1 2210
box -4 -6 84 206
use NAND3X1  _3144_
timestamp 1596033377
transform -1 0 1560 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3142_
timestamp 1596033377
transform 1 0 1560 0 -1 2210
box -4 -6 68 206
use FILL  SFILL14320x20100
timestamp 1596033377
transform -1 0 1448 0 -1 2210
box -4 -6 20 206
use FILL  SFILL14480x20100
timestamp 1596033377
transform -1 0 1464 0 -1 2210
box -4 -6 20 206
use FILL  SFILL14640x20100
timestamp 1596033377
transform -1 0 1480 0 -1 2210
box -4 -6 20 206
use FILL  SFILL14800x20100
timestamp 1596033377
transform -1 0 1496 0 -1 2210
box -4 -6 20 206
use AND2X2  _3113_
timestamp 1596033377
transform 1 0 1624 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3090_
timestamp 1596033377
transform -1 0 1752 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3168_
timestamp 1596033377
transform -1 0 1816 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3110_
timestamp 1596033377
transform -1 0 1880 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3114_
timestamp 1596033377
transform -1 0 1944 0 -1 2210
box -4 -6 68 206
use AOI22X1  _3169_
timestamp 1596033377
transform 1 0 1944 0 -1 2210
box -4 -6 84 206
use NAND3X1  _3170_
timestamp 1596033377
transform 1 0 2024 0 -1 2210
box -4 -6 68 206
use INVX1  _3424_
timestamp 1596033377
transform 1 0 2088 0 -1 2210
box -4 -6 36 206
use NAND3X1  _3120_
timestamp 1596033377
transform -1 0 2184 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3092_
timestamp 1596033377
transform 1 0 2184 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3167_
timestamp 1596033377
transform -1 0 2296 0 -1 2210
box -4 -6 52 206
use AND2X2  _2362_
timestamp 1596033377
transform -1 0 2360 0 -1 2210
box -4 -6 68 206
use XNOR2X1  _2417_
timestamp 1596033377
transform 1 0 2360 0 -1 2210
box -4 -6 116 206
use NAND2X1  _2419_
timestamp 1596033377
transform 1 0 2472 0 -1 2210
box -4 -6 52 206
use NOR2X1  _2391_
timestamp 1596033377
transform 1 0 2520 0 -1 2210
box -4 -6 52 206
use XOR2X1  _2371_
timestamp 1596033377
transform -1 0 2680 0 -1 2210
box -4 -6 116 206
use NOR2X1  _2373_
timestamp 1596033377
transform 1 0 2680 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3426_
timestamp 1596033377
transform -1 0 2776 0 -1 2210
box -4 -6 52 206
use XOR2X1  _2378_
timestamp 1596033377
transform 1 0 2776 0 -1 2210
box -4 -6 116 206
use XNOR2X1  _2406_
timestamp 1596033377
transform 1 0 2952 0 -1 2210
box -4 -6 116 206
use FILL  SFILL28880x20100
timestamp 1596033377
transform -1 0 2904 0 -1 2210
box -4 -6 20 206
use FILL  SFILL29040x20100
timestamp 1596033377
transform -1 0 2920 0 -1 2210
box -4 -6 20 206
use FILL  SFILL29200x20100
timestamp 1596033377
transform -1 0 2936 0 -1 2210
box -4 -6 20 206
use FILL  SFILL29360x20100
timestamp 1596033377
transform -1 0 2952 0 -1 2210
box -4 -6 20 206
use NAND2X1  _2407_
timestamp 1596033377
transform -1 0 3112 0 -1 2210
box -4 -6 52 206
use XNOR2X1  _2405_
timestamp 1596033377
transform -1 0 3224 0 -1 2210
box -4 -6 116 206
use BUFX2  BUFX2_insert97
timestamp 1596033377
transform -1 0 3272 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2121_
timestamp 1596033377
transform -1 0 3320 0 -1 2210
box -4 -6 52 206
use OAI21X1  _2122_
timestamp 1596033377
transform -1 0 3384 0 -1 2210
box -4 -6 68 206
use INVX1  _2120_
timestamp 1596033377
transform -1 0 3416 0 -1 2210
box -4 -6 36 206
use INVX1  _2132_
timestamp 1596033377
transform -1 0 3448 0 -1 2210
box -4 -6 36 206
use INVX1  _2123_
timestamp 1596033377
transform -1 0 3480 0 -1 2210
box -4 -6 36 206
use OAI21X1  _2125_
timestamp 1596033377
transform 1 0 3480 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert196
timestamp 1596033377
transform 1 0 3544 0 -1 2210
box -4 -6 52 206
use NAND2X1  _2136_
timestamp 1596033377
transform 1 0 3592 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert138
timestamp 1596033377
transform 1 0 3640 0 -1 2210
box -4 -6 52 206
use INVX1  _2117_
timestamp 1596033377
transform 1 0 3688 0 -1 2210
box -4 -6 36 206
use OAI21X1  _4604_
timestamp 1596033377
transform -1 0 3784 0 -1 2210
box -4 -6 68 206
use NAND2X1  _4588_
timestamp 1596033377
transform -1 0 3832 0 -1 2210
box -4 -6 52 206
use NAND2X1  _4594_
timestamp 1596033377
transform -1 0 3880 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert179
timestamp 1596033377
transform -1 0 3928 0 -1 2210
box -4 -6 52 206
use OAI21X1  _4595_
timestamp 1596033377
transform -1 0 3992 0 -1 2210
box -4 -6 68 206
use NAND3X1  _3537_
timestamp 1596033377
transform -1 0 4056 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3538_
timestamp 1596033377
transform -1 0 4104 0 -1 2210
box -4 -6 52 206
use AND2X2  _3558_
timestamp 1596033377
transform -1 0 4168 0 -1 2210
box -4 -6 68 206
use AND2X2  _3559_
timestamp 1596033377
transform 1 0 4168 0 -1 2210
box -4 -6 68 206
use AND2X2  _3556_
timestamp 1596033377
transform 1 0 4232 0 -1 2210
box -4 -6 68 206
use AND2X2  _3555_
timestamp 1596033377
transform -1 0 4360 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3454_
timestamp 1596033377
transform 1 0 4360 0 -1 2210
box -4 -6 52 206
use FILL  SFILL44080x20100
timestamp 1596033377
transform -1 0 4424 0 -1 2210
box -4 -6 20 206
use NOR2X1  _3544_
timestamp 1596033377
transform 1 0 4472 0 -1 2210
box -4 -6 52 206
use INVX1  _3543_
timestamp 1596033377
transform -1 0 4552 0 -1 2210
box -4 -6 36 206
use AND2X2  _3557_
timestamp 1596033377
transform -1 0 4616 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3504_
timestamp 1596033377
transform -1 0 4664 0 -1 2210
box -4 -6 52 206
use FILL  SFILL44240x20100
timestamp 1596033377
transform -1 0 4440 0 -1 2210
box -4 -6 20 206
use FILL  SFILL44400x20100
timestamp 1596033377
transform -1 0 4456 0 -1 2210
box -4 -6 20 206
use FILL  SFILL44560x20100
timestamp 1596033377
transform -1 0 4472 0 -1 2210
box -4 -6 20 206
use AND2X2  _3561_
timestamp 1596033377
transform -1 0 4728 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3510_
timestamp 1596033377
transform 1 0 4728 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4296_
timestamp 1596033377
transform 1 0 4776 0 -1 2210
box -4 -6 196 206
use NAND2X1  _3840_
timestamp 1596033377
transform 1 0 4968 0 -1 2210
box -4 -6 52 206
use OAI21X1  _3841_
timestamp 1596033377
transform -1 0 5080 0 -1 2210
box -4 -6 68 206
use AOI21X1  _3653_
timestamp 1596033377
transform 1 0 5080 0 -1 2210
box -4 -6 68 206
use NOR2X1  _3652_
timestamp 1596033377
transform -1 0 5192 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert10
timestamp 1596033377
transform -1 0 5240 0 -1 2210
box -4 -6 52 206
use MUX2X1  _3911_
timestamp 1596033377
transform 1 0 5240 0 -1 2210
box -4 -6 100 206
use MUX2X1  _4091_
timestamp 1596033377
transform 1 0 5336 0 -1 2210
box -4 -6 100 206
use BUFX2  BUFX2_insert273
timestamp 1596033377
transform 1 0 5432 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert69
timestamp 1596033377
transform -1 0 5528 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert68
timestamp 1596033377
transform -1 0 5576 0 -1 2210
box -4 -6 52 206
use NOR2X1  _3885_
timestamp 1596033377
transform -1 0 5624 0 -1 2210
box -4 -6 52 206
use AOI21X1  _3886_
timestamp 1596033377
transform -1 0 5688 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4334_
timestamp 1596033377
transform 1 0 5688 0 -1 2210
box -4 -6 196 206
use AND2X2  _3872_
timestamp 1596033377
transform -1 0 5944 0 -1 2210
box -4 -6 68 206
use NAND2X1  _3839_
timestamp 1596033377
transform 1 0 6008 0 -1 2210
box -4 -6 52 206
use FILL  SFILL59440x20100
timestamp 1596033377
transform -1 0 5960 0 -1 2210
box -4 -6 20 206
use FILL  SFILL59600x20100
timestamp 1596033377
transform -1 0 5976 0 -1 2210
box -4 -6 20 206
use FILL  SFILL59760x20100
timestamp 1596033377
transform -1 0 5992 0 -1 2210
box -4 -6 20 206
use FILL  SFILL59920x20100
timestamp 1596033377
transform -1 0 6008 0 -1 2210
box -4 -6 20 206
use AND2X2  _4263_
timestamp 1596033377
transform -1 0 6120 0 -1 2210
box -4 -6 68 206
use AND2X2  _3651_
timestamp 1596033377
transform 1 0 6120 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4318_
timestamp 1596033377
transform 1 0 6184 0 -1 2210
box -4 -6 196 206
use NOR2X1  _3703_
timestamp 1596033377
transform 1 0 6376 0 -1 2210
box -4 -6 52 206
use NAND2X1  _3751_
timestamp 1596033377
transform 1 0 6424 0 -1 2210
box -4 -6 52 206
use OAI21X1  _3752_
timestamp 1596033377
transform -1 0 6536 0 -1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert218
timestamp 1596033377
transform -1 0 6584 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert37
timestamp 1596033377
transform 1 0 6584 0 -1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert165
timestamp 1596033377
transform 1 0 6632 0 -1 2210
box -4 -6 52 206
use NOR2X1  _3808_
timestamp 1596033377
transform 1 0 6680 0 -1 2210
box -4 -6 52 206
use AOI21X1  _3809_
timestamp 1596033377
transform -1 0 6792 0 -1 2210
box -4 -6 68 206
use OAI21X1  _3708_
timestamp 1596033377
transform 1 0 6792 0 -1 2210
box -4 -6 68 206
use OAI21X1  _3709_
timestamp 1596033377
transform -1 0 6920 0 -1 2210
box -4 -6 68 206
use DFFPOSX1  _4361_
timestamp 1596033377
transform -1 0 7112 0 -1 2210
box -4 -6 196 206
use BUFX2  BUFX2_insert52
timestamp 1596033377
transform -1 0 7160 0 -1 2210
box -4 -6 52 206
use DFFPOSX1  _4376_
timestamp 1596033377
transform -1 0 7352 0 -1 2210
box -4 -6 196 206
use FILL  FILL70960x20100
timestamp 1596033377
transform -1 0 7368 0 -1 2210
box -4 -6 20 206
use FILL  FILL71120x20100
timestamp 1596033377
transform -1 0 7384 0 -1 2210
box -4 -6 20 206
use FILL  FILL71280x20100
timestamp 1596033377
transform -1 0 7400 0 -1 2210
box -4 -6 20 206
use NOR2X1  _3004_
timestamp 1596033377
transform 1 0 8 0 1 2210
box -4 -6 52 206
use INVX1  _2998_
timestamp 1596033377
transform -1 0 88 0 1 2210
box -4 -6 36 206
use OAI22X1  _3000_
timestamp 1596033377
transform 1 0 88 0 1 2210
box -4 -6 84 206
use INVX1  _2999_
timestamp 1596033377
transform -1 0 200 0 1 2210
box -4 -6 36 206
use INVX1  _3050_
timestamp 1596033377
transform 1 0 200 0 1 2210
box -4 -6 36 206
use OAI22X1  _3052_
timestamp 1596033377
transform 1 0 232 0 1 2210
box -4 -6 84 206
use INVX1  _3051_
timestamp 1596033377
transform -1 0 344 0 1 2210
box -4 -6 36 206
use NAND3X1  _3014_
timestamp 1596033377
transform 1 0 344 0 1 2210
box -4 -6 68 206
use AOI22X1  _3013_
timestamp 1596033377
transform -1 0 488 0 1 2210
box -4 -6 84 206
use NOR2X1  _3041_
timestamp 1596033377
transform 1 0 488 0 1 2210
box -4 -6 52 206
use NAND3X1  _3040_
timestamp 1596033377
transform 1 0 536 0 1 2210
box -4 -6 68 206
use AOI22X1  _3039_
timestamp 1596033377
transform -1 0 680 0 1 2210
box -4 -6 84 206
use AND2X2  _3035_
timestamp 1596033377
transform -1 0 744 0 1 2210
box -4 -6 68 206
use NAND3X1  _3034_
timestamp 1596033377
transform 1 0 744 0 1 2210
box -4 -6 68 206
use NAND3X1  _3008_
timestamp 1596033377
transform 1 0 808 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert64
timestamp 1596033377
transform -1 0 920 0 1 2210
box -4 -6 52 206
use AND2X2  _2973_
timestamp 1596033377
transform -1 0 984 0 1 2210
box -4 -6 68 206
use NAND3X1  _3042_
timestamp 1596033377
transform -1 0 1048 0 1 2210
box -4 -6 68 206
use BUFX2  BUFX2_insert234
timestamp 1596033377
transform -1 0 1096 0 1 2210
box -4 -6 52 206
use INVX1  _3442_
timestamp 1596033377
transform 1 0 1096 0 1 2210
box -4 -6 36 206
use AND2X2  _2968_
timestamp 1596033377
transform -1 0 1192 0 1 2210
box -4 -6 68 206
use NOR2X1  _2960_
timestamp 1596033377
transform 1 0 1192 0 1 2210
box -4 -6 52 206
use AND2X2  _2972_
timestamp 1596033377
transform -1 0 1304 0 1 2210
box -4 -6 68 206
use NOR2X1  _2975_
timestamp 1596033377
transform -1 0 1352 0 1 2210
box -4 -6 52 206
use XOR2X1  _2290_
timestamp 1596033377
transform -1 0 1464 0 1 2210
box -4 -6 116 206
use NAND3X1  _2977_
timestamp 1596033377
transform -1 0 1592 0 1 2210
box -4 -6 68 206
use NAND3X1  _2980_
timestamp 1596033377
transform -1 0 1656 0 1 2210
box -4 -6 68 206
use FILL  SFILL14640x22100
timestamp 1596033377
transform 1 0 1464 0 1 2210
box -4 -6 20 206
use FILL  SFILL14800x22100
timestamp 1596033377
transform 1 0 1480 0 1 2210
box -4 -6 20 206
use FILL  SFILL14960x22100
timestamp 1596033377
transform 1 0 1496 0 1 2210
box -4 -6 20 206
use FILL  SFILL15120x22100
timestamp 1596033377
transform 1 0 1512 0 1 2210
box -4 -6 20 206
use NAND2X1  _2974_
timestamp 1596033377
transform -1 0 1704 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert224
timestamp 1596033377
transform -1 0 1752 0 1 2210
box -4 -6 52 206
use OR2X2  _2339_
timestamp 1596033377
transform 1 0 1752 0 1 2210
box -4 -6 68 206
use INVX1  _2939_
timestamp 1596033377
transform 1 0 1816 0 1 2210
box -4 -6 36 206
use OAI22X1  _2950_
timestamp 1596033377
transform 1 0 1848 0 1 2210
box -4 -6 84 206
use INVX1  _2940_
timestamp 1596033377
transform -1 0 1960 0 1 2210
box -4 -6 36 206
use NAND2X1  _3109_
timestamp 1596033377
transform -1 0 2008 0 1 2210
box -4 -6 52 206
use NAND3X1  _3116_
timestamp 1596033377
transform -1 0 2072 0 1 2210
box -4 -6 68 206
use NOR2X1  _3119_
timestamp 1596033377
transform 1 0 2072 0 1 2210
box -4 -6 52 206
use NAND3X1  _3118_
timestamp 1596033377
transform 1 0 2120 0 1 2210
box -4 -6 68 206
use AOI22X1  _3091_
timestamp 1596033377
transform -1 0 2264 0 1 2210
box -4 -6 84 206
use NAND2X1  _3089_
timestamp 1596033377
transform -1 0 2312 0 1 2210
box -4 -6 52 206
use INVX1  _3076_
timestamp 1596033377
transform 1 0 2312 0 1 2210
box -4 -6 36 206
use NOR2X1  _3082_
timestamp 1596033377
transform -1 0 2392 0 1 2210
box -4 -6 52 206
use OAI22X1  _3078_
timestamp 1596033377
transform 1 0 2392 0 1 2210
box -4 -6 84 206
use INVX1  _3077_
timestamp 1596033377
transform 1 0 2472 0 1 2210
box -4 -6 36 206
use AND2X2  _2359_
timestamp 1596033377
transform -1 0 2568 0 1 2210
box -4 -6 68 206
use XOR2X1  _2389_
timestamp 1596033377
transform 1 0 2568 0 1 2210
box -4 -6 116 206
use OR2X2  _3425_
timestamp 1596033377
transform 1 0 2680 0 1 2210
box -4 -6 68 206
use OAI21X1  _3443_
timestamp 1596033377
transform -1 0 2808 0 1 2210
box -4 -6 68 206
use XOR2X1  _2377_
timestamp 1596033377
transform 1 0 2808 0 1 2210
box -4 -6 116 206
use OAI21X1  _3499_
timestamp 1596033377
transform -1 0 3048 0 1 2210
box -4 -6 68 206
use FILL  SFILL29200x22100
timestamp 1596033377
transform 1 0 2920 0 1 2210
box -4 -6 20 206
use FILL  SFILL29360x22100
timestamp 1596033377
transform 1 0 2936 0 1 2210
box -4 -6 20 206
use FILL  SFILL29520x22100
timestamp 1596033377
transform 1 0 2952 0 1 2210
box -4 -6 20 206
use FILL  SFILL29680x22100
timestamp 1596033377
transform 1 0 2968 0 1 2210
box -4 -6 20 206
use OAI21X1  _3534_
timestamp 1596033377
transform -1 0 3112 0 1 2210
box -4 -6 68 206
use OAI21X1  _3506_
timestamp 1596033377
transform -1 0 3176 0 1 2210
box -4 -6 68 206
use OAI21X1  _3527_
timestamp 1596033377
transform 1 0 3176 0 1 2210
box -4 -6 68 206
use OAI21X1  _3520_
timestamp 1596033377
transform -1 0 3304 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4427_
timestamp 1596033377
transform -1 0 3496 0 1 2210
box -4 -6 196 206
use NAND2X1  _2124_
timestamp 1596033377
transform 1 0 3496 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert293
timestamp 1596033377
transform 1 0 3544 0 1 2210
box -4 -6 52 206
use NAND3X1  _4474_
timestamp 1596033377
transform -1 0 3656 0 1 2210
box -4 -6 68 206
use OAI21X1  _4129_
timestamp 1596033377
transform 1 0 3656 0 1 2210
box -4 -6 68 206
use AOI21X1  _4130_
timestamp 1596033377
transform -1 0 3784 0 1 2210
box -4 -6 68 206
use OAI21X1  _4589_
timestamp 1596033377
transform -1 0 3848 0 1 2210
box -4 -6 68 206
use NAND2X1  _4591_
timestamp 1596033377
transform -1 0 3896 0 1 2210
box -4 -6 52 206
use OAI21X1  _4592_
timestamp 1596033377
transform -1 0 3960 0 1 2210
box -4 -6 68 206
use NAND3X1  _3530_
timestamp 1596033377
transform -1 0 4024 0 1 2210
box -4 -6 68 206
use INVX1  _4590_
timestamp 1596033377
transform -1 0 4056 0 1 2210
box -4 -6 36 206
use INVX1  _4587_
timestamp 1596033377
transform -1 0 4088 0 1 2210
box -4 -6 36 206
use INVX1  _4614_
timestamp 1596033377
transform -1 0 4120 0 1 2210
box -4 -6 36 206
use NAND2X1  _3532_
timestamp 1596033377
transform -1 0 4168 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert128
timestamp 1596033377
transform 1 0 4168 0 1 2210
box -4 -6 52 206
use NAND2X1  _3448_
timestamp 1596033377
transform 1 0 4216 0 1 2210
box -4 -6 52 206
use INVX1  _4626_
timestamp 1596033377
transform 1 0 4264 0 1 2210
box -4 -6 36 206
use NOR2X1  _3546_
timestamp 1596033377
transform 1 0 4296 0 1 2210
box -4 -6 52 206
use INVX1  _3545_
timestamp 1596033377
transform -1 0 4376 0 1 2210
box -4 -6 36 206
use NAND3X1  _3523_
timestamp 1596033377
transform -1 0 4440 0 1 2210
box -4 -6 68 206
use INVX4  _3660_
timestamp 1596033377
transform 1 0 4504 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert127
timestamp 1596033377
transform 1 0 4552 0 1 2210
box -4 -6 52 206
use NAND3X1  _3446_
timestamp 1596033377
transform -1 0 4664 0 1 2210
box -4 -6 68 206
use FILL  SFILL44400x22100
timestamp 1596033377
transform 1 0 4440 0 1 2210
box -4 -6 20 206
use FILL  SFILL44560x22100
timestamp 1596033377
transform 1 0 4456 0 1 2210
box -4 -6 20 206
use FILL  SFILL44720x22100
timestamp 1596033377
transform 1 0 4472 0 1 2210
box -4 -6 20 206
use FILL  SFILL44880x22100
timestamp 1596033377
transform 1 0 4488 0 1 2210
box -4 -6 20 206
use NAND3X1  _3502_
timestamp 1596033377
transform -1 0 4728 0 1 2210
box -4 -6 68 206
use MUX2X1  _3928_
timestamp 1596033377
transform -1 0 4824 0 1 2210
box -4 -6 100 206
use DFFPOSX1  _4392_
timestamp 1596033377
transform -1 0 5016 0 1 2210
box -4 -6 196 206
use NOR2X1  _3925_
timestamp 1596033377
transform 1 0 5016 0 1 2210
box -4 -6 52 206
use OAI22X1  _3927_
timestamp 1596033377
transform 1 0 5064 0 1 2210
box -4 -6 84 206
use OAI21X1  _3926_
timestamp 1596033377
transform -1 0 5208 0 1 2210
box -4 -6 68 206
use MUX2X1  _3924_
timestamp 1596033377
transform -1 0 5304 0 1 2210
box -4 -6 100 206
use MUX2X1  _4102_
timestamp 1596033377
transform -1 0 5400 0 1 2210
box -4 -6 100 206
use NOR2X1  _4103_
timestamp 1596033377
transform 1 0 5400 0 1 2210
box -4 -6 52 206
use OAI22X1  _4105_
timestamp 1596033377
transform 1 0 5448 0 1 2210
box -4 -6 84 206
use OAI21X1  _4104_
timestamp 1596033377
transform -1 0 5592 0 1 2210
box -4 -6 68 206
use MUX2X1  _4106_
timestamp 1596033377
transform -1 0 5688 0 1 2210
box -4 -6 100 206
use NOR2X1  _3875_
timestamp 1596033377
transform 1 0 5688 0 1 2210
box -4 -6 52 206
use AOI21X1  _3876_
timestamp 1596033377
transform -1 0 5800 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4329_
timestamp 1596033377
transform -1 0 5992 0 1 2210
box -4 -6 196 206
use FILL  SFILL59920x22100
timestamp 1596033377
transform 1 0 5992 0 1 2210
box -4 -6 20 206
use FILL  SFILL60080x22100
timestamp 1596033377
transform 1 0 6008 0 1 2210
box -4 -6 20 206
use BUFX2  BUFX2_insert206
timestamp 1596033377
transform -1 0 6104 0 1 2210
box -4 -6 52 206
use BUFX2  BUFX2_insert118
timestamp 1596033377
transform 1 0 6104 0 1 2210
box -4 -6 52 206
use OAI22X1  _4101_
timestamp 1596033377
transform -1 0 6232 0 1 2210
box -4 -6 84 206
use FILL  SFILL60240x22100
timestamp 1596033377
transform 1 0 6024 0 1 2210
box -4 -6 20 206
use FILL  SFILL60400x22100
timestamp 1596033377
transform 1 0 6040 0 1 2210
box -4 -6 20 206
use NOR2X1  _4099_
timestamp 1596033377
transform 1 0 6232 0 1 2210
box -4 -6 52 206
use OAI21X1  _4100_
timestamp 1596033377
transform -1 0 6344 0 1 2210
box -4 -6 68 206
use MUX2X1  _4098_
timestamp 1596033377
transform 1 0 6344 0 1 2210
box -4 -6 100 206
use OAI21X1  _3922_
timestamp 1596033377
transform 1 0 6440 0 1 2210
box -4 -6 68 206
use OAI22X1  _3923_
timestamp 1596033377
transform 1 0 6504 0 1 2210
box -4 -6 84 206
use NOR2X1  _3921_
timestamp 1596033377
transform 1 0 6584 0 1 2210
box -4 -6 52 206
use MUX2X1  _3920_
timestamp 1596033377
transform 1 0 6632 0 1 2210
box -4 -6 100 206
use DFFPOSX1  _4377_
timestamp 1596033377
transform -1 0 6920 0 1 2210
box -4 -6 196 206
use OAI21X1  _3718_
timestamp 1596033377
transform 1 0 6920 0 1 2210
box -4 -6 68 206
use DFFPOSX1  _4366_
timestamp 1596033377
transform -1 0 7176 0 1 2210
box -4 -6 196 206
use DFFPOSX1  _4408_
timestamp 1596033377
transform -1 0 7368 0 1 2210
box -4 -6 196 206
use FILL  FILL71120x22100
timestamp 1596033377
transform 1 0 7368 0 1 2210
box -4 -6 20 206
use FILL  FILL71280x22100
timestamp 1596033377
transform 1 0 7384 0 1 2210
box -4 -6 20 206
use INVX1  _3001_
timestamp 1596033377
transform 1 0 8 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3003_
timestamp 1596033377
transform 1 0 40 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3002_
timestamp 1596033377
transform -1 0 152 0 -1 2610
box -4 -6 52 206
use INVX1  _3053_
timestamp 1596033377
transform 1 0 152 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3055_
timestamp 1596033377
transform 1 0 184 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3054_
timestamp 1596033377
transform -1 0 296 0 -1 2610
box -4 -6 52 206
use NAND3X1  _3064_
timestamp 1596033377
transform 1 0 296 0 -1 2610
box -4 -6 68 206
use NAND3X1  _3012_
timestamp 1596033377
transform 1 0 360 0 -1 2610
box -4 -6 68 206
use NAND3X1  _3038_
timestamp 1596033377
transform -1 0 488 0 -1 2610
box -4 -6 68 206
use INVX1  _3027_
timestamp 1596033377
transform 1 0 488 0 -1 2610
box -4 -6 36 206
use OAI21X1  _3029_
timestamp 1596033377
transform 1 0 520 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3028_
timestamp 1596033377
transform -1 0 632 0 -1 2610
box -4 -6 52 206
use NOR2X1  _3030_
timestamp 1596033377
transform -1 0 680 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert114
timestamp 1596033377
transform -1 0 728 0 -1 2610
box -4 -6 52 206
use NAND3X1  _3060_
timestamp 1596033377
transform -1 0 792 0 -1 2610
box -4 -6 68 206
use NAND3X1  _3372_
timestamp 1596033377
transform -1 0 856 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3132_
timestamp 1596033377
transform 1 0 856 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3133_
timestamp 1596033377
transform -1 0 968 0 -1 2610
box -4 -6 68 206
use INVX1  _3131_
timestamp 1596033377
transform -1 0 1000 0 -1 2610
box -4 -6 36 206
use BUFX2  BUFX2_insert215
timestamp 1596033377
transform -1 0 1048 0 -1 2610
box -4 -6 52 206
use NOR2X1  _3134_
timestamp 1596033377
transform -1 0 1096 0 -1 2610
box -4 -6 52 206
use INVX1  _3129_
timestamp 1596033377
transform 1 0 1096 0 -1 2610
box -4 -6 36 206
use OAI22X1  _3130_
timestamp 1596033377
transform -1 0 1208 0 -1 2610
box -4 -6 84 206
use INVX1  _3128_
timestamp 1596033377
transform -1 0 1240 0 -1 2610
box -4 -6 36 206
use INVX1  _3498_
timestamp 1596033377
transform 1 0 1240 0 -1 2610
box -4 -6 36 206
use NAND2X1  _2981_
timestamp 1596033377
transform 1 0 1272 0 -1 2610
box -4 -6 52 206
use NOR3X1  _2985_
timestamp 1596033377
transform -1 0 1448 0 -1 2610
box -4 -6 132 206
use NAND2X1  _2942_
timestamp 1596033377
transform -1 0 1560 0 -1 2610
box -4 -6 52 206
use INVX1  _2941_
timestamp 1596033377
transform -1 0 1592 0 -1 2610
box -4 -6 36 206
use NOR2X1  _2953_
timestamp 1596033377
transform -1 0 1640 0 -1 2610
box -4 -6 52 206
use FILL  SFILL14480x24100
timestamp 1596033377
transform -1 0 1464 0 -1 2610
box -4 -6 20 206
use FILL  SFILL14640x24100
timestamp 1596033377
transform -1 0 1480 0 -1 2610
box -4 -6 20 206
use FILL  SFILL14800x24100
timestamp 1596033377
transform -1 0 1496 0 -1 2610
box -4 -6 20 206
use FILL  SFILL14960x24100
timestamp 1596033377
transform -1 0 1512 0 -1 2610
box -4 -6 20 206
use BUFX2  BUFX2_insert113
timestamp 1596033377
transform 1 0 1640 0 -1 2610
box -4 -6 52 206
use AND2X2  _2355_
timestamp 1596033377
transform -1 0 1752 0 -1 2610
box -4 -6 68 206
use XOR2X1  _2433_
timestamp 1596033377
transform 1 0 1752 0 -1 2610
box -4 -6 116 206
use INVX1  _2951_
timestamp 1596033377
transform 1 0 1864 0 -1 2610
box -4 -6 36 206
use NOR2X1  _2957_
timestamp 1596033377
transform -1 0 1944 0 -1 2610
box -4 -6 52 206
use OAI22X1  _2956_
timestamp 1596033377
transform 1 0 1944 0 -1 2610
box -4 -6 84 206
use NAND3X1  _2990_
timestamp 1596033377
transform 1 0 2024 0 -1 2610
box -4 -6 68 206
use NOR2X1  _3108_
timestamp 1596033377
transform 1 0 2088 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3107_
timestamp 1596033377
transform -1 0 2200 0 -1 2610
box -4 -6 68 206
use NAND2X1  _2965_
timestamp 1596033377
transform -1 0 2248 0 -1 2610
box -4 -6 52 206
use AOI22X1  _3117_
timestamp 1596033377
transform -1 0 2328 0 -1 2610
box -4 -6 84 206
use OAI21X1  _3081_
timestamp 1596033377
transform -1 0 2392 0 -1 2610
box -4 -6 68 206
use INVX1  _3079_
timestamp 1596033377
transform -1 0 2424 0 -1 2610
box -4 -6 36 206
use NOR2X1  _3160_
timestamp 1596033377
transform 1 0 2424 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3159_
timestamp 1596033377
transform -1 0 2536 0 -1 2610
box -4 -6 68 206
use INVX1  _3157_
timestamp 1596033377
transform -1 0 2568 0 -1 2610
box -4 -6 36 206
use XNOR2X1  _2428_
timestamp 1596033377
transform 1 0 2568 0 -1 2610
box -4 -6 116 206
use XNOR2X1  _2429_
timestamp 1596033377
transform -1 0 2792 0 -1 2610
box -4 -6 116 206
use NOR3X1  _2384_
timestamp 1596033377
transform 1 0 2792 0 -1 2610
box -4 -6 132 206
use INVX1  _3533_
timestamp 1596033377
transform 1 0 2984 0 -1 2610
box -4 -6 36 206
use FILL  SFILL29200x24100
timestamp 1596033377
transform -1 0 2936 0 -1 2610
box -4 -6 20 206
use FILL  SFILL29360x24100
timestamp 1596033377
transform -1 0 2952 0 -1 2610
box -4 -6 20 206
use FILL  SFILL29520x24100
timestamp 1596033377
transform -1 0 2968 0 -1 2610
box -4 -6 20 206
use FILL  SFILL29680x24100
timestamp 1596033377
transform -1 0 2984 0 -1 2610
box -4 -6 20 206
use NOR3X1  _2416_
timestamp 1596033377
transform -1 0 3144 0 -1 2610
box -4 -6 132 206
use INVX1  _3519_
timestamp 1596033377
transform 1 0 3144 0 -1 2610
box -4 -6 36 206
use DFFPOSX1  _4568_
timestamp 1596033377
transform 1 0 3176 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  _4567_
timestamp 1596033377
transform -1 0 3560 0 -1 2610
box -4 -6 196 206
use AOI21X1  _4477_
timestamp 1596033377
transform -1 0 3624 0 -1 2610
box -4 -6 68 206
use INVX1  _4472_
timestamp 1596033377
transform 1 0 3624 0 -1 2610
box -4 -6 36 206
use AOI22X1  _4476_
timestamp 1596033377
transform -1 0 3736 0 -1 2610
box -4 -6 84 206
use NAND3X1  _4475_
timestamp 1596033377
transform 1 0 3736 0 -1 2610
box -4 -6 68 206
use AOI22X1  _4483_
timestamp 1596033377
transform -1 0 3880 0 -1 2610
box -4 -6 84 206
use OAI21X1  _4473_
timestamp 1596033377
transform -1 0 3944 0 -1 2610
box -4 -6 68 206
use NAND2X1  _4467_
timestamp 1596033377
transform -1 0 3992 0 -1 2610
box -4 -6 52 206
use INVX1  _4466_
timestamp 1596033377
transform -1 0 4024 0 -1 2610
box -4 -6 36 206
use INVX1  _4457_
timestamp 1596033377
transform -1 0 4056 0 -1 2610
box -4 -6 36 206
use NAND2X1  _4460_
timestamp 1596033377
transform 1 0 4056 0 -1 2610
box -4 -6 52 206
use AOI21X1  _4465_
timestamp 1596033377
transform -1 0 4168 0 -1 2610
box -4 -6 68 206
use AOI22X1  _4464_
timestamp 1596033377
transform -1 0 4248 0 -1 2610
box -4 -6 84 206
use DFFPOSX1  _4566_
timestamp 1596033377
transform -1 0 4440 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_insert180
timestamp 1596033377
transform 1 0 4504 0 -1 2610
box -4 -6 52 206
use NAND3X1  _3516_
timestamp 1596033377
transform -1 0 4616 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3517_
timestamp 1596033377
transform -1 0 4664 0 -1 2610
box -4 -6 52 206
use FILL  SFILL44400x24100
timestamp 1596033377
transform -1 0 4456 0 -1 2610
box -4 -6 20 206
use FILL  SFILL44560x24100
timestamp 1596033377
transform -1 0 4472 0 -1 2610
box -4 -6 20 206
use FILL  SFILL44720x24100
timestamp 1596033377
transform -1 0 4488 0 -1 2610
box -4 -6 20 206
use FILL  SFILL44880x24100
timestamp 1596033377
transform -1 0 4504 0 -1 2610
box -4 -6 20 206
use NAND2X1  _3511_
timestamp 1596033377
transform -1 0 4712 0 -1 2610
box -4 -6 52 206
use AND2X2  _3560_
timestamp 1596033377
transform 1 0 4712 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3483_
timestamp 1596033377
transform -1 0 4824 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3524_
timestamp 1596033377
transform 1 0 4824 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3503_
timestamp 1596033377
transform 1 0 4872 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3531_
timestamp 1596033377
transform -1 0 4968 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3525_
timestamp 1596033377
transform -1 0 5016 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3441_
timestamp 1596033377
transform 1 0 5016 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3447_
timestamp 1596033377
transform 1 0 5064 0 -1 2610
box -4 -6 52 206
use INVX4  _3657_
timestamp 1596033377
transform 1 0 5112 0 -1 2610
box -4 -6 52 206
use NAND2X1  _3842_
timestamp 1596033377
transform -1 0 5208 0 -1 2610
box -4 -6 52 206
use MUX2X1  _3950_
timestamp 1596033377
transform -1 0 5304 0 -1 2610
box -4 -6 100 206
use MUX2X1  _4128_
timestamp 1596033377
transform -1 0 5400 0 -1 2610
box -4 -6 100 206
use AOI21X1  _3656_
timestamp 1596033377
transform 1 0 5400 0 -1 2610
box -4 -6 68 206
use NOR2X1  _3655_
timestamp 1596033377
transform 1 0 5464 0 -1 2610
box -4 -6 52 206
use AOI21X1  _4267_
timestamp 1596033377
transform -1 0 5576 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4409_
timestamp 1596033377
transform -1 0 5768 0 -1 2610
box -4 -6 196 206
use BUFX2  BUFX2_insert219
timestamp 1596033377
transform -1 0 5816 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert163
timestamp 1596033377
transform 1 0 5816 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert278
timestamp 1596033377
transform -1 0 5912 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert256
timestamp 1596033377
transform 1 0 5976 0 -1 2610
box -4 -6 52 206
use FILL  SFILL59120x24100
timestamp 1596033377
transform -1 0 5928 0 -1 2610
box -4 -6 20 206
use FILL  SFILL59280x24100
timestamp 1596033377
transform -1 0 5944 0 -1 2610
box -4 -6 20 206
use FILL  SFILL59440x24100
timestamp 1596033377
transform -1 0 5960 0 -1 2610
box -4 -6 20 206
use FILL  SFILL59600x24100
timestamp 1596033377
transform -1 0 5976 0 -1 2610
box -4 -6 20 206
use NOR2X1  _4268_
timestamp 1596033377
transform -1 0 6072 0 -1 2610
box -4 -6 52 206
use AOI21X1  _4269_
timestamp 1596033377
transform -1 0 6136 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4410_
timestamp 1596033377
transform -1 0 6328 0 -1 2610
box -4 -6 196 206
use NOR2X1  _3943_
timestamp 1596033377
transform 1 0 6328 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert143
timestamp 1596033377
transform 1 0 6376 0 -1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert258
timestamp 1596033377
transform 1 0 6424 0 -1 2610
box -4 -6 52 206
use OAI22X1  _3945_
timestamp 1596033377
transform 1 0 6472 0 -1 2610
box -4 -6 84 206
use OAI21X1  _3944_
timestamp 1596033377
transform -1 0 6616 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4315_
timestamp 1596033377
transform -1 0 6808 0 -1 2610
box -4 -6 196 206
use OAI21X1  _3746_
timestamp 1596033377
transform -1 0 6872 0 -1 2610
box -4 -6 68 206
use NAND2X1  _3741_
timestamp 1596033377
transform 1 0 6872 0 -1 2610
box -4 -6 52 206
use OAI21X1  _3742_
timestamp 1596033377
transform -1 0 6984 0 -1 2610
box -4 -6 68 206
use DFFPOSX1  _4313_
timestamp 1596033377
transform -1 0 7176 0 -1 2610
box -4 -6 196 206
use DFFPOSX1  _4345_
timestamp 1596033377
transform -1 0 7368 0 -1 2610
box -4 -6 196 206
use FILL  FILL71120x24100
timestamp 1596033377
transform -1 0 7384 0 -1 2610
box -4 -6 20 206
use FILL  FILL71280x24100
timestamp 1596033377
transform -1 0 7400 0 -1 2610
box -4 -6 20 206
use INVX1  _3313_
timestamp 1596033377
transform 1 0 8 0 1 2610
box -4 -6 36 206
use OAI21X1  _3315_
timestamp 1596033377
transform 1 0 40 0 1 2610
box -4 -6 68 206
use NAND2X1  _3314_
timestamp 1596033377
transform -1 0 152 0 1 2610
box -4 -6 52 206
use INVX1  _3310_
timestamp 1596033377
transform 1 0 152 0 1 2610
box -4 -6 36 206
use OAI22X1  _3312_
timestamp 1596033377
transform 1 0 184 0 1 2610
box -4 -6 84 206
use INVX1  _3311_
timestamp 1596033377
transform -1 0 296 0 1 2610
box -4 -6 36 206
use NOR2X1  _3316_
timestamp 1596033377
transform -1 0 344 0 1 2610
box -4 -6 52 206
use AOI22X1  _3247_
timestamp 1596033377
transform 1 0 344 0 1 2610
box -4 -6 84 206
use NAND3X1  _3248_
timestamp 1596033377
transform -1 0 488 0 1 2610
box -4 -6 68 206
use NAND3X1  _3246_
timestamp 1596033377
transform 1 0 488 0 1 2610
box -4 -6 68 206
use NAND3X1  _3328_
timestamp 1596033377
transform 1 0 552 0 1 2610
box -4 -6 68 206
use INVX1  _3024_
timestamp 1596033377
transform 1 0 616 0 1 2610
box -4 -6 36 206
use OAI22X1  _3026_
timestamp 1596033377
transform 1 0 648 0 1 2610
box -4 -6 84 206
use INVX1  _3025_
timestamp 1596033377
transform -1 0 760 0 1 2610
box -4 -6 36 206
use NAND3X1  _3376_
timestamp 1596033377
transform 1 0 760 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert112
timestamp 1596033377
transform 1 0 824 0 1 2610
box -4 -6 52 206
use NAND2X1  _2949_
timestamp 1596033377
transform 1 0 872 0 1 2610
box -4 -6 52 206
use NAND2X1  _2955_
timestamp 1596033377
transform 1 0 920 0 1 2610
box -4 -6 52 206
use NAND2X1  _2954_
timestamp 1596033377
transform 1 0 968 0 1 2610
box -4 -6 52 206
use NAND2X1  _2947_
timestamp 1596033377
transform 1 0 1016 0 1 2610
box -4 -6 52 206
use NAND2X1  _2961_
timestamp 1596033377
transform -1 0 1112 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert271
timestamp 1596033377
transform -1 0 1160 0 1 2610
box -4 -6 52 206
use INVX1  _2946_
timestamp 1596033377
transform -1 0 1192 0 1 2610
box -4 -6 36 206
use NOR2X1  _2948_
timestamp 1596033377
transform 1 0 1192 0 1 2610
box -4 -6 52 206
use NAND2X1  _2945_
timestamp 1596033377
transform -1 0 1288 0 1 2610
box -4 -6 52 206
use INVX1  _2944_
timestamp 1596033377
transform -1 0 1320 0 1 2610
box -4 -6 36 206
use INVX8  _2943_
timestamp 1596033377
transform -1 0 1400 0 1 2610
box -4 -6 84 206
use FILL  SFILL14000x26100
timestamp 1596033377
transform 1 0 1400 0 1 2610
box -4 -6 20 206
use NOR2X1  _2982_
timestamp 1596033377
transform 1 0 1464 0 1 2610
box -4 -6 52 206
use BUFX2  BUFX2_insert111
timestamp 1596033377
transform -1 0 1560 0 1 2610
box -4 -6 52 206
use AND2X2  _2979_
timestamp 1596033377
transform -1 0 1624 0 1 2610
box -4 -6 68 206
use FILL  SFILL14160x26100
timestamp 1596033377
transform 1 0 1416 0 1 2610
box -4 -6 20 206
use FILL  SFILL14320x26100
timestamp 1596033377
transform 1 0 1432 0 1 2610
box -4 -6 20 206
use FILL  SFILL14480x26100
timestamp 1596033377
transform 1 0 1448 0 1 2610
box -4 -6 20 206
use NOR2X1  _2989_
timestamp 1596033377
transform 1 0 1624 0 1 2610
box -4 -6 52 206
use NAND2X1  _2983_
timestamp 1596033377
transform 1 0 1672 0 1 2610
box -4 -6 52 206
use NAND3X1  _2988_
timestamp 1596033377
transform -1 0 1784 0 1 2610
box -4 -6 68 206
use NOR2X1  _2966_
timestamp 1596033377
transform -1 0 1832 0 1 2610
box -4 -6 52 206
use NOR3X1  _2986_
timestamp 1596033377
transform 1 0 1832 0 1 2610
box -4 -6 132 206
use INVX1  _3102_
timestamp 1596033377
transform 1 0 1960 0 1 2610
box -4 -6 36 206
use OAI22X1  _3104_
timestamp 1596033377
transform 1 0 1992 0 1 2610
box -4 -6 84 206
use INVX1  _3103_
timestamp 1596033377
transform -1 0 2104 0 1 2610
box -4 -6 36 206
use NAND2X1  _3106_
timestamp 1596033377
transform 1 0 2104 0 1 2610
box -4 -6 52 206
use INVX1  _3105_
timestamp 1596033377
transform 1 0 2152 0 1 2610
box -4 -6 36 206
use NAND2X1  _3080_
timestamp 1596033377
transform 1 0 2184 0 1 2610
box -4 -6 52 206
use INVX1  _3155_
timestamp 1596033377
transform 1 0 2232 0 1 2610
box -4 -6 36 206
use OAI22X1  _3156_
timestamp 1596033377
transform -1 0 2344 0 1 2610
box -4 -6 84 206
use INVX1  _3154_
timestamp 1596033377
transform -1 0 2376 0 1 2610
box -4 -6 36 206
use INVX1  _2952_
timestamp 1596033377
transform -1 0 2408 0 1 2610
box -4 -6 36 206
use NAND2X1  _3158_
timestamp 1596033377
transform 1 0 2408 0 1 2610
box -4 -6 52 206
use NAND2X1  _2432_
timestamp 1596033377
transform -1 0 2504 0 1 2610
box -4 -6 52 206
use NOR3X1  _2431_
timestamp 1596033377
transform 1 0 2504 0 1 2610
box -4 -6 132 206
use NAND3X1  _2430_
timestamp 1596033377
transform 1 0 2632 0 1 2610
box -4 -6 68 206
use NAND3X1  _2385_
timestamp 1596033377
transform 1 0 2696 0 1 2610
box -4 -6 68 206
use OAI21X1  _3492_
timestamp 1596033377
transform 1 0 2760 0 1 2610
box -4 -6 68 206
use OAI21X1  _3485_
timestamp 1596033377
transform -1 0 2888 0 1 2610
box -4 -6 68 206
use OAI21X1  _3513_
timestamp 1596033377
transform 1 0 2888 0 1 2610
box -4 -6 68 206
use FILL  SFILL29520x26100
timestamp 1596033377
transform 1 0 2952 0 1 2610
box -4 -6 20 206
use FILL  SFILL29680x26100
timestamp 1596033377
transform 1 0 2968 0 1 2610
box -4 -6 20 206
use FILL  SFILL29840x26100
timestamp 1596033377
transform 1 0 2984 0 1 2610
box -4 -6 20 206
use FILL  SFILL30000x26100
timestamp 1596033377
transform 1 0 3000 0 1 2610
box -4 -6 20 206
use DFFPOSX1  _4571_
timestamp 1596033377
transform 1 0 3016 0 1 2610
box -4 -6 196 206
use AOI21X1  _4504_
timestamp 1596033377
transform -1 0 3272 0 1 2610
box -4 -6 68 206
use AOI21X1  _4484_
timestamp 1596033377
transform -1 0 3336 0 1 2610
box -4 -6 68 206
use NAND3X1  _4482_
timestamp 1596033377
transform 1 0 3336 0 1 2610
box -4 -6 68 206
use AOI22X1  _4503_
timestamp 1596033377
transform -1 0 3480 0 1 2610
box -4 -6 84 206
use INVX2  _4478_
timestamp 1596033377
transform 1 0 3480 0 1 2610
box -4 -6 36 206
use INVX1  _4481_
timestamp 1596033377
transform -1 0 3544 0 1 2610
box -4 -6 36 206
use NOR2X1  _4480_
timestamp 1596033377
transform 1 0 3544 0 1 2610
box -4 -6 52 206
use OAI21X1  _4479_
timestamp 1596033377
transform -1 0 3656 0 1 2610
box -4 -6 68 206
use NAND2X1  _4468_
timestamp 1596033377
transform 1 0 3656 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _4565_
timestamp 1596033377
transform -1 0 3896 0 1 2610
box -4 -6 196 206
use NAND3X1  _4469_
timestamp 1596033377
transform 1 0 3896 0 1 2610
box -4 -6 68 206
use AOI21X1  _4471_
timestamp 1596033377
transform 1 0 3960 0 1 2610
box -4 -6 68 206
use AOI22X1  _4470_
timestamp 1596033377
transform -1 0 4104 0 1 2610
box -4 -6 84 206
use INVX1  _4605_
timestamp 1596033377
transform -1 0 4136 0 1 2610
box -4 -6 36 206
use NAND3X1  _3488_
timestamp 1596033377
transform -1 0 4200 0 1 2610
box -4 -6 68 206
use NAND2X1  _4627_
timestamp 1596033377
transform -1 0 4248 0 1 2610
box -4 -6 52 206
use OAI21X1  _4628_
timestamp 1596033377
transform -1 0 4312 0 1 2610
box -4 -6 68 206
use NAND3X1  _3495_
timestamp 1596033377
transform -1 0 4376 0 1 2610
box -4 -6 68 206
use INVX1  _4623_
timestamp 1596033377
transform -1 0 4408 0 1 2610
box -4 -6 36 206
use FILL  SFILL44080x26100
timestamp 1596033377
transform 1 0 4408 0 1 2610
box -4 -6 20 206
use INVX4  _3687_
timestamp 1596033377
transform -1 0 4520 0 1 2610
box -4 -6 52 206
use INVX1  _4617_
timestamp 1596033377
transform 1 0 4520 0 1 2610
box -4 -6 36 206
use NAND2X1  _3497_
timestamp 1596033377
transform -1 0 4600 0 1 2610
box -4 -6 52 206
use INVX4  _3693_
timestamp 1596033377
transform -1 0 4648 0 1 2610
box -4 -6 52 206
use FILL  SFILL44240x26100
timestamp 1596033377
transform 1 0 4424 0 1 2610
box -4 -6 20 206
use FILL  SFILL44400x26100
timestamp 1596033377
transform 1 0 4440 0 1 2610
box -4 -6 20 206
use FILL  SFILL44560x26100
timestamp 1596033377
transform 1 0 4456 0 1 2610
box -4 -6 20 206
use NAND2X1  _3489_
timestamp 1596033377
transform -1 0 4696 0 1 2610
box -4 -6 52 206
use NAND2X1  _3518_
timestamp 1596033377
transform 1 0 4696 0 1 2610
box -4 -6 52 206
use CLKBUF1  CLKBUF1_insert30
timestamp 1596033377
transform 1 0 4744 0 1 2610
box -4 -6 148 206
use INVX4  _3684_
timestamp 1596033377
transform -1 0 4936 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _4297_
timestamp 1596033377
transform -1 0 5128 0 1 2610
box -4 -6 196 206
use OAI21X1  _3843_
timestamp 1596033377
transform 1 0 5128 0 1 2610
box -4 -6 68 206
use BUFX2  BUFX2_insert9
timestamp 1596033377
transform -1 0 5240 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _4393_
timestamp 1596033377
transform -1 0 5432 0 1 2610
box -4 -6 196 206
use NOR2X1  _4266_
timestamp 1596033377
transform -1 0 5480 0 1 2610
box -4 -6 52 206
use AOI21X1  _3659_
timestamp 1596033377
transform 1 0 5480 0 1 2610
box -4 -6 68 206
use NOR2X1  _3658_
timestamp 1596033377
transform -1 0 5592 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _4394_
timestamp 1596033377
transform 1 0 5592 0 1 2610
box -4 -6 196 206
use MUX2X1  _4117_
timestamp 1596033377
transform -1 0 5880 0 1 2610
box -4 -6 100 206
use MUX2X1  _4113_
timestamp 1596033377
transform 1 0 5880 0 1 2610
box -4 -6 100 206
use FILL  SFILL59760x26100
timestamp 1596033377
transform 1 0 5976 0 1 2610
box -4 -6 20 206
use FILL  SFILL59920x26100
timestamp 1596033377
transform 1 0 5992 0 1 2610
box -4 -6 20 206
use FILL  SFILL60080x26100
timestamp 1596033377
transform 1 0 6008 0 1 2610
box -4 -6 20 206
use MUX2X1  _3935_
timestamp 1596033377
transform -1 0 6136 0 1 2610
box -4 -6 100 206
use BUFX2  BUFX2_insert89
timestamp 1596033377
transform 1 0 6136 0 1 2610
box -4 -6 52 206
use OAI22X1  _4123_
timestamp 1596033377
transform -1 0 6264 0 1 2610
box -4 -6 84 206
use FILL  SFILL60240x26100
timestamp 1596033377
transform 1 0 6024 0 1 2610
box -4 -6 20 206
use NOR2X1  _4121_
timestamp 1596033377
transform -1 0 6312 0 1 2610
box -4 -6 52 206
use OAI21X1  _4122_
timestamp 1596033377
transform -1 0 6376 0 1 2610
box -4 -6 68 206
use OAI22X1  _4112_
timestamp 1596033377
transform -1 0 6456 0 1 2610
box -4 -6 84 206
use NOR2X1  _4110_
timestamp 1596033377
transform -1 0 6504 0 1 2610
box -4 -6 52 206
use OAI21X1  _3710_
timestamp 1596033377
transform 1 0 6504 0 1 2610
box -4 -6 68 206
use OAI21X1  _3711_
timestamp 1596033377
transform -1 0 6632 0 1 2610
box -4 -6 68 206
use NAND2X1  _3745_
timestamp 1596033377
transform 1 0 6632 0 1 2610
box -4 -6 52 206
use DFFPOSX1  _4362_
timestamp 1596033377
transform -1 0 6872 0 1 2610
box -4 -6 196 206
use OAI21X1  _3712_
timestamp 1596033377
transform 1 0 6872 0 1 2610
box -4 -6 68 206
use OAI21X1  _3713_
timestamp 1596033377
transform -1 0 7000 0 1 2610
box -4 -6 68 206
use DFFPOSX1  _4363_
timestamp 1596033377
transform -1 0 7192 0 1 2610
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert22
timestamp 1596033377
transform -1 0 7336 0 1 2610
box -4 -6 148 206
use NAND2X1  _3775_
timestamp 1596033377
transform -1 0 7384 0 1 2610
box -4 -6 52 206
use FILL  FILL71280x26100
timestamp 1596033377
transform 1 0 7384 0 1 2610
box -4 -6 20 206
use INVX1  _3365_
timestamp 1596033377
transform 1 0 8 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3367_
timestamp 1596033377
transform 1 0 40 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3366_
timestamp 1596033377
transform -1 0 152 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3368_
timestamp 1596033377
transform -1 0 200 0 -1 3010
box -4 -6 52 206
use INVX1  _3362_
timestamp 1596033377
transform 1 0 200 0 -1 3010
box -4 -6 36 206
use OAI22X1  _3364_
timestamp 1596033377
transform 1 0 232 0 -1 3010
box -4 -6 84 206
use INVX1  _3363_
timestamp 1596033377
transform -1 0 344 0 -1 3010
box -4 -6 36 206
use NAND3X1  _3250_
timestamp 1596033377
transform 1 0 344 0 -1 3010
box -4 -6 68 206
use NOR2X1  _3249_
timestamp 1596033377
transform 1 0 408 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3380_
timestamp 1596033377
transform 1 0 456 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3377_
timestamp 1596033377
transform 1 0 520 0 -1 3010
box -4 -6 84 206
use NOR2X1  _3379_
timestamp 1596033377
transform -1 0 648 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3378_
timestamp 1596033377
transform -1 0 712 0 -1 3010
box -4 -6 68 206
use INVX1  _3287_
timestamp 1596033377
transform 1 0 712 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3289_
timestamp 1596033377
transform 1 0 744 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3288_
timestamp 1596033377
transform -1 0 856 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3290_
timestamp 1596033377
transform -1 0 904 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert226
timestamp 1596033377
transform -1 0 952 0 -1 3010
box -4 -6 52 206
use INVX1  _3285_
timestamp 1596033377
transform 1 0 952 0 -1 3010
box -4 -6 36 206
use OAI22X1  _3286_
timestamp 1596033377
transform -1 0 1064 0 -1 3010
box -4 -6 84 206
use INVX1  _3284_
timestamp 1596033377
transform -1 0 1096 0 -1 3010
box -4 -6 36 206
use NAND2X1  _2962_
timestamp 1596033377
transform -1 0 1144 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert237
timestamp 1596033377
transform 1 0 1144 0 -1 3010
box -4 -6 52 206
use NAND2X1  _2969_
timestamp 1596033377
transform -1 0 1240 0 -1 3010
box -4 -6 52 206
use NAND3X1  _3320_
timestamp 1596033377
transform 1 0 1240 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3317_
timestamp 1596033377
transform 1 0 1304 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert65
timestamp 1596033377
transform -1 0 1400 0 -1 3010
box -4 -6 52 206
use FILL  SFILL14000x28100
timestamp 1596033377
transform -1 0 1416 0 -1 3010
box -4 -6 20 206
use BUFX2  BUFX2_insert236
timestamp 1596033377
transform 1 0 1464 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert63
timestamp 1596033377
transform -1 0 1560 0 -1 3010
box -4 -6 52 206
use NAND2X1  _2826_
timestamp 1596033377
transform 1 0 1560 0 -1 3010
box -4 -6 52 206
use AOI22X1  _2844_
timestamp 1596033377
transform -1 0 1688 0 -1 3010
box -4 -6 84 206
use FILL  SFILL14160x28100
timestamp 1596033377
transform -1 0 1432 0 -1 3010
box -4 -6 20 206
use FILL  SFILL14320x28100
timestamp 1596033377
transform -1 0 1448 0 -1 3010
box -4 -6 20 206
use FILL  SFILL14480x28100
timestamp 1596033377
transform -1 0 1464 0 -1 3010
box -4 -6 20 206
use AOI22X1  _2987_
timestamp 1596033377
transform 1 0 1688 0 -1 3010
box -4 -6 84 206
use NAND3X1  _2978_
timestamp 1596033377
transform -1 0 1832 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3187_
timestamp 1596033377
transform 1 0 1832 0 -1 3010
box -4 -6 52 206
use INVX1  _2964_
timestamp 1596033377
transform 1 0 1880 0 -1 3010
box -4 -6 36 206
use NAND3X1  _2984_
timestamp 1596033377
transform -1 0 1976 0 -1 3010
box -4 -6 68 206
use AOI22X1  _3221_
timestamp 1596033377
transform 1 0 1976 0 -1 3010
box -4 -6 84 206
use AOI22X1  _3351_
timestamp 1596033377
transform 1 0 2056 0 -1 3010
box -4 -6 84 206
use OAI21X1  _2970_
timestamp 1596033377
transform 1 0 2136 0 -1 3010
box -4 -6 68 206
use NOR2X1  _2971_
timestamp 1596033377
transform -1 0 2248 0 -1 3010
box -4 -6 52 206
use INVX1  _2959_
timestamp 1596033377
transform -1 0 2280 0 -1 3010
box -4 -6 36 206
use OAI22X1  _2963_
timestamp 1596033377
transform -1 0 2360 0 -1 3010
box -4 -6 84 206
use INVX1  _2958_
timestamp 1596033377
transform -1 0 2392 0 -1 3010
box -4 -6 36 206
use NAND2X1  _2967_
timestamp 1596033377
transform -1 0 2440 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3184_
timestamp 1596033377
transform 1 0 2440 0 -1 3010
box -4 -6 52 206
use INVX1  _3181_
timestamp 1596033377
transform 1 0 2488 0 -1 3010
box -4 -6 36 206
use OAI22X1  _3182_
timestamp 1596033377
transform -1 0 2600 0 -1 3010
box -4 -6 84 206
use INVX1  _3180_
timestamp 1596033377
transform -1 0 2632 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3262_
timestamp 1596033377
transform 1 0 2632 0 -1 3010
box -4 -6 52 206
use NAND2X1  _3210_
timestamp 1596033377
transform -1 0 2728 0 -1 3010
box -4 -6 52 206
use NOR2X1  _2401_
timestamp 1596033377
transform 1 0 2728 0 -1 3010
box -4 -6 52 206
use INVX1  _3491_
timestamp 1596033377
transform 1 0 2776 0 -1 3010
box -4 -6 36 206
use INVX1  _3484_
timestamp 1596033377
transform 1 0 2808 0 -1 3010
box -4 -6 36 206
use OAI21X1  _3211_
timestamp 1596033377
transform -1 0 2904 0 -1 3010
box -4 -6 68 206
use INVX1  _3512_
timestamp 1596033377
transform 1 0 2904 0 -1 3010
box -4 -6 36 206
use INVX1  _3209_
timestamp 1596033377
transform -1 0 3032 0 -1 3010
box -4 -6 36 206
use FILL  SFILL29360x28100
timestamp 1596033377
transform -1 0 2952 0 -1 3010
box -4 -6 20 206
use FILL  SFILL29520x28100
timestamp 1596033377
transform -1 0 2968 0 -1 3010
box -4 -6 20 206
use FILL  SFILL29680x28100
timestamp 1596033377
transform -1 0 2984 0 -1 3010
box -4 -6 20 206
use FILL  SFILL29840x28100
timestamp 1596033377
transform -1 0 3000 0 -1 3010
box -4 -6 20 206
use NAND3X1  _2415_
timestamp 1596033377
transform -1 0 3096 0 -1 3010
box -4 -6 68 206
use INVX1  _3505_
timestamp 1596033377
transform 1 0 3096 0 -1 3010
box -4 -6 36 206
use INVX1  _3526_
timestamp 1596033377
transform 1 0 3128 0 -1 3010
box -4 -6 36 206
use NAND3X1  _4502_
timestamp 1596033377
transform -1 0 3224 0 -1 3010
box -4 -6 68 206
use OAI21X1  _4500_
timestamp 1596033377
transform -1 0 3288 0 -1 3010
box -4 -6 68 206
use NOR3X1  _4514_
timestamp 1596033377
transform -1 0 3416 0 -1 3010
box -4 -6 132 206
use INVX1  _4499_
timestamp 1596033377
transform 1 0 3416 0 -1 3010
box -4 -6 36 206
use INVX1  _4492_
timestamp 1596033377
transform -1 0 3480 0 -1 3010
box -4 -6 36 206
use AOI21X1  _4498_
timestamp 1596033377
transform -1 0 3544 0 -1 3010
box -4 -6 68 206
use NAND3X1  _4496_
timestamp 1596033377
transform 1 0 3544 0 -1 3010
box -4 -6 68 206
use OAI21X1  _4493_
timestamp 1596033377
transform -1 0 3672 0 -1 3010
box -4 -6 68 206
use AOI22X1  _4497_
timestamp 1596033377
transform -1 0 3752 0 -1 3010
box -4 -6 84 206
use NOR3X1  _4494_
timestamp 1596033377
transform 1 0 3752 0 -1 3010
box -4 -6 132 206
use NAND3X1  _4488_
timestamp 1596033377
transform 1 0 3880 0 -1 3010
box -4 -6 68 206
use INVX1  _4487_
timestamp 1596033377
transform -1 0 3976 0 -1 3010
box -4 -6 36 206
use OAI21X1  _4486_
timestamp 1596033377
transform 1 0 3976 0 -1 3010
box -4 -6 68 206
use NAND3X1  _4489_
timestamp 1596033377
transform -1 0 4104 0 -1 3010
box -4 -6 68 206
use AOI21X1  _4491_
timestamp 1596033377
transform 1 0 4104 0 -1 3010
box -4 -6 68 206
use AOI22X1  _4490_
timestamp 1596033377
transform -1 0 4248 0 -1 3010
box -4 -6 84 206
use INVX1  _4461_
timestamp 1596033377
transform -1 0 4280 0 -1 3010
box -4 -6 36 206
use NOR2X1  _4459_
timestamp 1596033377
transform 1 0 4280 0 -1 3010
box -4 -6 52 206
use NOR2X1  _4463_
timestamp 1596033377
transform -1 0 4376 0 -1 3010
box -4 -6 52 206
use NAND2X1  _4558_
timestamp 1596033377
transform -1 0 4424 0 -1 3010
box -4 -6 52 206
use INVX1  _4458_
timestamp 1596033377
transform -1 0 4520 0 -1 3010
box -4 -6 36 206
use INVX4  _4456_
timestamp 1596033377
transform 1 0 4520 0 -1 3010
box -4 -6 52 206
use INVX1  _4608_
timestamp 1596033377
transform -1 0 4600 0 -1 3010
box -4 -6 36 206
use NAND2X1  _3496_
timestamp 1596033377
transform -1 0 4648 0 -1 3010
box -4 -6 52 206
use FILL  SFILL44240x28100
timestamp 1596033377
transform -1 0 4440 0 -1 3010
box -4 -6 20 206
use FILL  SFILL44400x28100
timestamp 1596033377
transform -1 0 4456 0 -1 3010
box -4 -6 20 206
use FILL  SFILL44560x28100
timestamp 1596033377
transform -1 0 4472 0 -1 3010
box -4 -6 20 206
use FILL  SFILL44720x28100
timestamp 1596033377
transform -1 0 4488 0 -1 3010
box -4 -6 20 206
use NAND2X1  _3490_
timestamp 1596033377
transform -1 0 4696 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4395_
timestamp 1596033377
transform 1 0 4696 0 -1 3010
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert25
timestamp 1596033377
transform -1 0 5032 0 -1 3010
box -4 -6 148 206
use DFFPOSX1  _4411_
timestamp 1596033377
transform 1 0 5032 0 -1 3010
box -4 -6 196 206
use AOI21X1  _4271_
timestamp 1596033377
transform 1 0 5224 0 -1 3010
box -4 -6 68 206
use NOR2X1  _4270_
timestamp 1596033377
transform 1 0 5288 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3847_
timestamp 1596033377
transform 1 0 5336 0 -1 3010
box -4 -6 68 206
use NAND2X1  _3846_
timestamp 1596033377
transform -1 0 5448 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4299_
timestamp 1596033377
transform 1 0 5448 0 -1 3010
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert28
timestamp 1596033377
transform 1 0 5640 0 -1 3010
box -4 -6 148 206
use BUFX2  BUFX2_insert164
timestamp 1596033377
transform -1 0 5832 0 -1 3010
box -4 -6 52 206
use NOR2X1  _3879_
timestamp 1596033377
transform -1 0 5880 0 -1 3010
box -4 -6 52 206
use OAI21X1  _4126_
timestamp 1596033377
transform 1 0 5880 0 -1 3010
box -4 -6 68 206
use OAI22X1  _4116_
timestamp 1596033377
transform -1 0 6088 0 -1 3010
box -4 -6 84 206
use FILL  SFILL59440x28100
timestamp 1596033377
transform -1 0 5960 0 -1 3010
box -4 -6 20 206
use FILL  SFILL59600x28100
timestamp 1596033377
transform -1 0 5976 0 -1 3010
box -4 -6 20 206
use FILL  SFILL59760x28100
timestamp 1596033377
transform -1 0 5992 0 -1 3010
box -4 -6 20 206
use FILL  SFILL59920x28100
timestamp 1596033377
transform -1 0 6008 0 -1 3010
box -4 -6 20 206
use INVX8  _4087_
timestamp 1596033377
transform -1 0 6168 0 -1 3010
box -4 -6 84 206
use BUFX2  BUFX2_insert117
timestamp 1596033377
transform 1 0 6168 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert207
timestamp 1596033377
transform 1 0 6216 0 -1 3010
box -4 -6 52 206
use MUX2X1  _3939_
timestamp 1596033377
transform -1 0 6360 0 -1 3010
box -4 -6 100 206
use OAI21X1  _4115_
timestamp 1596033377
transform -1 0 6424 0 -1 3010
box -4 -6 68 206
use OAI21X1  _4111_
timestamp 1596033377
transform -1 0 6488 0 -1 3010
box -4 -6 68 206
use MUX2X1  _3942_
timestamp 1596033377
transform -1 0 6584 0 -1 3010
box -4 -6 100 206
use MUX2X1  _4120_
timestamp 1596033377
transform -1 0 6680 0 -1 3010
box -4 -6 100 206
use MUX2X1  _4109_
timestamp 1596033377
transform 1 0 6680 0 -1 3010
box -4 -6 100 206
use DFFPOSX1  _4346_
timestamp 1596033377
transform -1 0 6968 0 -1 3010
box -4 -6 196 206
use NAND2X1  _3777_
timestamp 1596033377
transform 1 0 6968 0 -1 3010
box -4 -6 52 206
use OAI21X1  _3778_
timestamp 1596033377
transform -1 0 7080 0 -1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert4
timestamp 1596033377
transform -1 0 7128 0 -1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert8
timestamp 1596033377
transform 1 0 7128 0 -1 3010
box -4 -6 52 206
use DFFPOSX1  _4347_
timestamp 1596033377
transform -1 0 7368 0 -1 3010
box -4 -6 196 206
use FILL  FILL71120x28100
timestamp 1596033377
transform -1 0 7384 0 -1 3010
box -4 -6 20 206
use FILL  FILL71280x28100
timestamp 1596033377
transform -1 0 7400 0 -1 3010
box -4 -6 20 206
use INVX1  _3235_
timestamp 1596033377
transform 1 0 8 0 1 3010
box -4 -6 36 206
use OAI21X1  _3237_
timestamp 1596033377
transform 1 0 40 0 1 3010
box -4 -6 68 206
use NAND2X1  _3236_
timestamp 1596033377
transform -1 0 152 0 1 3010
box -4 -6 52 206
use INVX1  _3359_
timestamp 1596033377
transform 1 0 152 0 1 3010
box -4 -6 36 206
use OAI22X1  _3360_
timestamp 1596033377
transform -1 0 264 0 1 3010
box -4 -6 84 206
use NOR2X1  _3238_
timestamp 1596033377
transform -1 0 312 0 1 3010
box -4 -6 52 206
use INVX1  _3233_
timestamp 1596033377
transform 1 0 312 0 1 3010
box -4 -6 36 206
use OAI22X1  _3234_
timestamp 1596033377
transform -1 0 424 0 1 3010
box -4 -6 84 206
use INVX1  _3232_
timestamp 1596033377
transform -1 0 456 0 1 3010
box -4 -6 36 206
use NOR2X1  _3361_
timestamp 1596033377
transform 1 0 456 0 1 3010
box -4 -6 52 206
use INVX1  _3356_
timestamp 1596033377
transform 1 0 504 0 1 3010
box -4 -6 36 206
use OAI22X1  _3357_
timestamp 1596033377
transform -1 0 616 0 1 3010
box -4 -6 84 206
use INVX1  _3355_
timestamp 1596033377
transform 1 0 616 0 1 3010
box -4 -6 36 206
use NAND2X1  _3245_
timestamp 1596033377
transform 1 0 648 0 1 3010
box -4 -6 52 206
use NOR2X1  _3327_
timestamp 1596033377
transform -1 0 744 0 1 3010
box -4 -6 52 206
use NAND2X1  _3375_
timestamp 1596033377
transform -1 0 792 0 1 3010
box -4 -6 52 206
use NAND3X1  _3298_
timestamp 1596033377
transform 1 0 792 0 1 3010
box -4 -6 68 206
use NAND3X1  _3324_
timestamp 1596033377
transform 1 0 856 0 1 3010
box -4 -6 68 206
use AOI22X1  _3325_
timestamp 1596033377
transform -1 0 1000 0 1 3010
box -4 -6 84 206
use AOI22X1  _3299_
timestamp 1596033377
transform -1 0 1080 0 1 3010
box -4 -6 84 206
use NAND2X1  _3369_
timestamp 1596033377
transform 1 0 1080 0 1 3010
box -4 -6 52 206
use NAND3X1  _3374_
timestamp 1596033377
transform 1 0 1128 0 1 3010
box -4 -6 68 206
use AND2X2  _3373_
timestamp 1596033377
transform 1 0 1192 0 1 3010
box -4 -6 68 206
use AND2X2  _3321_
timestamp 1596033377
transform 1 0 1256 0 1 3010
box -4 -6 68 206
use NAND3X1  _3322_
timestamp 1596033377
transform 1 0 1320 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert227
timestamp 1596033377
transform -1 0 1432 0 1 3010
box -4 -6 52 206
use NAND3X1  _3242_
timestamp 1596033377
transform 1 0 1496 0 1 3010
box -4 -6 68 206
use NAND3X1  _3294_
timestamp 1596033377
transform 1 0 1560 0 1 3010
box -4 -6 68 206
use FILL  SFILL14320x30100
timestamp 1596033377
transform 1 0 1432 0 1 3010
box -4 -6 20 206
use FILL  SFILL14480x30100
timestamp 1596033377
transform 1 0 1448 0 1 3010
box -4 -6 20 206
use FILL  SFILL14640x30100
timestamp 1596033377
transform 1 0 1464 0 1 3010
box -4 -6 20 206
use FILL  SFILL14800x30100
timestamp 1596033377
transform 1 0 1480 0 1 3010
box -4 -6 20 206
use NAND3X1  _3268_
timestamp 1596033377
transform 1 0 1624 0 1 3010
box -4 -6 68 206
use NAND3X1  _3190_
timestamp 1596033377
transform 1 0 1688 0 1 3010
box -4 -6 68 206
use NAND3X1  _3216_
timestamp 1596033377
transform 1 0 1752 0 1 3010
box -4 -6 68 206
use NAND3X1  _3346_
timestamp 1596033377
transform 1 0 1816 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert223
timestamp 1596033377
transform 1 0 1880 0 1 3010
box -4 -6 52 206
use NAND3X1  _3272_
timestamp 1596033377
transform 1 0 1928 0 1 3010
box -4 -6 68 206
use AOI22X1  _3273_
timestamp 1596033377
transform -1 0 2072 0 1 3010
box -4 -6 84 206
use NAND3X1  _3220_
timestamp 1596033377
transform 1 0 2072 0 1 3010
box -4 -6 68 206
use NAND3X1  _3352_
timestamp 1596033377
transform -1 0 2200 0 1 3010
box -4 -6 68 206
use NAND3X1  _3350_
timestamp 1596033377
transform -1 0 2264 0 1 3010
box -4 -6 68 206
use NAND3X1  _3194_
timestamp 1596033377
transform -1 0 2328 0 1 3010
box -4 -6 68 206
use AOI22X1  _3195_
timestamp 1596033377
transform 1 0 2328 0 1 3010
box -4 -6 84 206
use NAND3X1  _3196_
timestamp 1596033377
transform 1 0 2408 0 1 3010
box -4 -6 68 206
use NOR2X1  _3197_
timestamp 1596033377
transform -1 0 2520 0 1 3010
box -4 -6 52 206
use NAND3X1  _3198_
timestamp 1596033377
transform 1 0 2520 0 1 3010
box -4 -6 68 206
use NOR2X1  _3186_
timestamp 1596033377
transform 1 0 2584 0 1 3010
box -4 -6 52 206
use OAI21X1  _3185_
timestamp 1596033377
transform -1 0 2696 0 1 3010
box -4 -6 68 206
use INVX1  _3183_
timestamp 1596033377
transform -1 0 2728 0 1 3010
box -4 -6 36 206
use NAND3X1  _2400_
timestamp 1596033377
transform -1 0 2792 0 1 3010
box -4 -6 68 206
use OAI21X1  _3263_
timestamp 1596033377
transform -1 0 2856 0 1 3010
box -4 -6 68 206
use INVX1  _3261_
timestamp 1596033377
transform -1 0 2888 0 1 3010
box -4 -6 36 206
use NOR2X1  _3212_
timestamp 1596033377
transform -1 0 2936 0 1 3010
box -4 -6 52 206
use OAI22X1  _3208_
timestamp 1596033377
transform 1 0 3000 0 1 3010
box -4 -6 84 206
use FILL  SFILL29360x30100
timestamp 1596033377
transform 1 0 2936 0 1 3010
box -4 -6 20 206
use FILL  SFILL29520x30100
timestamp 1596033377
transform 1 0 2952 0 1 3010
box -4 -6 20 206
use FILL  SFILL29680x30100
timestamp 1596033377
transform 1 0 2968 0 1 3010
box -4 -6 20 206
use FILL  SFILL29840x30100
timestamp 1596033377
transform 1 0 2984 0 1 3010
box -4 -6 20 206
use INVX1  _3207_
timestamp 1596033377
transform 1 0 3080 0 1 3010
box -4 -6 36 206
use XNOR2X1  _2408_
timestamp 1596033377
transform 1 0 3112 0 1 3010
box -4 -6 116 206
use DFFPOSX1  _4570_
timestamp 1596033377
transform 1 0 3224 0 1 3010
box -4 -6 196 206
use AOI21X1  _4511_
timestamp 1596033377
transform -1 0 3480 0 1 3010
box -4 -6 68 206
use NAND3X1  _4509_
timestamp 1596033377
transform -1 0 3544 0 1 3010
box -4 -6 68 206
use OAI21X1  _4506_
timestamp 1596033377
transform -1 0 3608 0 1 3010
box -4 -6 68 206
use NAND3X1  _4501_
timestamp 1596033377
transform 1 0 3608 0 1 3010
box -4 -6 68 206
use NAND2X1  _4495_
timestamp 1596033377
transform 1 0 3672 0 1 3010
box -4 -6 52 206
use AOI22X1  _4510_
timestamp 1596033377
transform -1 0 3800 0 1 3010
box -4 -6 84 206
use INVX1  _2126_
timestamp 1596033377
transform -1 0 3832 0 1 3010
box -4 -6 36 206
use INVX1  _4485_
timestamp 1596033377
transform -1 0 3864 0 1 3010
box -4 -6 36 206
use DFFPOSX1  _4569_
timestamp 1596033377
transform -1 0 4056 0 1 3010
box -4 -6 196 206
use INVX1  _4611_
timestamp 1596033377
transform -1 0 4088 0 1 3010
box -4 -6 36 206
use INVX1  _4559_
timestamp 1596033377
transform 1 0 4088 0 1 3010
box -4 -6 36 206
use OAI21X1  _4560_
timestamp 1596033377
transform -1 0 4184 0 1 3010
box -4 -6 68 206
use NAND3X1  _4562_
timestamp 1596033377
transform -1 0 4248 0 1 3010
box -4 -6 68 206
use NAND3X1  _4563_
timestamp 1596033377
transform -1 0 4312 0 1 3010
box -4 -6 68 206
use NOR2X1  _4462_
timestamp 1596033377
transform -1 0 4360 0 1 3010
box -4 -6 52 206
use AOI21X1  _4564_
timestamp 1596033377
transform 1 0 4360 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4580_
timestamp 1596033377
transform -1 0 4680 0 1 3010
box -4 -6 196 206
use FILL  SFILL44240x30100
timestamp 1596033377
transform 1 0 4424 0 1 3010
box -4 -6 20 206
use FILL  SFILL44400x30100
timestamp 1596033377
transform 1 0 4440 0 1 3010
box -4 -6 20 206
use FILL  SFILL44560x30100
timestamp 1596033377
transform 1 0 4456 0 1 3010
box -4 -6 20 206
use FILL  SFILL44720x30100
timestamp 1596033377
transform 1 0 4472 0 1 3010
box -4 -6 20 206
use INVX1  _4620_
timestamp 1596033377
transform -1 0 4712 0 1 3010
box -4 -6 36 206
use AOI21X1  _3662_
timestamp 1596033377
transform 1 0 4712 0 1 3010
box -4 -6 68 206
use NOR2X1  _3661_
timestamp 1596033377
transform -1 0 4824 0 1 3010
box -4 -6 52 206
use INVX4  _3690_
timestamp 1596033377
transform -1 0 4872 0 1 3010
box -4 -6 52 206
use DFFPOSX1  _4298_
timestamp 1596033377
transform 1 0 4872 0 1 3010
box -4 -6 196 206
use OAI21X1  _3845_
timestamp 1596033377
transform -1 0 5128 0 1 3010
box -4 -6 68 206
use NAND2X1  _3844_
timestamp 1596033377
transform -1 0 5176 0 1 3010
box -4 -6 52 206
use MUX2X1  _3946_
timestamp 1596033377
transform 1 0 5176 0 1 3010
box -4 -6 100 206
use MUX2X1  _4124_
timestamp 1596033377
transform -1 0 5368 0 1 3010
box -4 -6 100 206
use OAI22X1  _4127_
timestamp 1596033377
transform -1 0 5448 0 1 3010
box -4 -6 84 206
use NOR2X1  _4125_
timestamp 1596033377
transform -1 0 5496 0 1 3010
box -4 -6 52 206
use OAI22X1  _3949_
timestamp 1596033377
transform -1 0 5576 0 1 3010
box -4 -6 84 206
use NOR2X1  _3947_
timestamp 1596033377
transform 1 0 5576 0 1 3010
box -4 -6 52 206
use INVX4  _3675_
timestamp 1596033377
transform 1 0 5624 0 1 3010
box -4 -6 52 206
use BUFX2  BUFX2_insert11
timestamp 1596033377
transform -1 0 5720 0 1 3010
box -4 -6 52 206
use OAI21X1  _3948_
timestamp 1596033377
transform -1 0 5784 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4331_
timestamp 1596033377
transform -1 0 5976 0 1 3010
box -4 -6 196 206
use FILL  SFILL59760x30100
timestamp 1596033377
transform 1 0 5976 0 1 3010
box -4 -6 20 206
use FILL  SFILL59920x30100
timestamp 1596033377
transform 1 0 5992 0 1 3010
box -4 -6 20 206
use FILL  SFILL60080x30100
timestamp 1596033377
transform 1 0 6008 0 1 3010
box -4 -6 20 206
use NOR2X1  _4114_
timestamp 1596033377
transform -1 0 6088 0 1 3010
box -4 -6 52 206
use AOI21X1  _3880_
timestamp 1596033377
transform -1 0 6152 0 1 3010
box -4 -6 68 206
use BUFX2  BUFX2_insert71
timestamp 1596033377
transform -1 0 6200 0 1 3010
box -4 -6 52 206
use NOR2X1  _3936_
timestamp 1596033377
transform 1 0 6200 0 1 3010
box -4 -6 52 206
use FILL  SFILL60240x30100
timestamp 1596033377
transform 1 0 6024 0 1 3010
box -4 -6 20 206
use OAI22X1  _3938_
timestamp 1596033377
transform 1 0 6248 0 1 3010
box -4 -6 84 206
use OAI21X1  _3937_
timestamp 1596033377
transform -1 0 6392 0 1 3010
box -4 -6 68 206
use INVX8  _3907_
timestamp 1596033377
transform -1 0 6472 0 1 3010
box -4 -6 84 206
use NOR2X1  _3932_
timestamp 1596033377
transform -1 0 6520 0 1 3010
box -4 -6 52 206
use OAI22X1  _3934_
timestamp 1596033377
transform 1 0 6520 0 1 3010
box -4 -6 84 206
use OAI21X1  _3933_
timestamp 1596033377
transform -1 0 6664 0 1 3010
box -4 -6 68 206
use NOR2X1  _3812_
timestamp 1596033377
transform 1 0 6664 0 1 3010
box -4 -6 52 206
use AOI21X1  _3813_
timestamp 1596033377
transform -1 0 6776 0 1 3010
box -4 -6 68 206
use MUX2X1  _3931_
timestamp 1596033377
transform -1 0 6872 0 1 3010
box -4 -6 100 206
use NAND2X1  _3743_
timestamp 1596033377
transform -1 0 6920 0 1 3010
box -4 -6 52 206
use OAI21X1  _3744_
timestamp 1596033377
transform -1 0 6984 0 1 3010
box -4 -6 68 206
use AOI21X1  _4293_
timestamp 1596033377
transform -1 0 7048 0 1 3010
box -4 -6 68 206
use DFFPOSX1  _4314_
timestamp 1596033377
transform -1 0 7240 0 1 3010
box -4 -6 196 206
use AOI21X1  _3878_
timestamp 1596033377
transform 1 0 7240 0 1 3010
box -4 -6 68 206
use NOR2X1  _3832_
timestamp 1596033377
transform -1 0 7352 0 1 3010
box -4 -6 52 206
use NOR2X1  _3877_
timestamp 1596033377
transform -1 0 7400 0 1 3010
box -4 -6 52 206
use INVX1  _3226_
timestamp 1596033377
transform 1 0 8 0 -1 3410
box -4 -6 36 206
use INVX1  _3358_
timestamp 1596033377
transform 1 0 40 0 -1 3410
box -4 -6 36 206
use NOR2X1  _3231_
timestamp 1596033377
transform 1 0 72 0 -1 3410
box -4 -6 52 206
use OAI22X1  _3227_
timestamp 1596033377
transform -1 0 200 0 -1 3410
box -4 -6 84 206
use INVX1  _3225_
timestamp 1596033377
transform -1 0 232 0 -1 3410
box -4 -6 36 206
use OR2X2  _2349_
timestamp 1596033377
transform -1 0 296 0 -1 3410
box -4 -6 68 206
use NOR2X1  _2321_
timestamp 1596033377
transform 1 0 296 0 -1 3410
box -4 -6 52 206
use NOR2X1  _2323_
timestamp 1596033377
transform 1 0 344 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3240_
timestamp 1596033377
transform 1 0 392 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3244_
timestamp 1596033377
transform 1 0 456 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3309_
timestamp 1596033377
transform 1 0 520 0 -1 3410
box -4 -6 52 206
use INVX1  _3304_
timestamp 1596033377
transform 1 0 568 0 -1 3410
box -4 -6 36 206
use OAI22X1  _3305_
timestamp 1596033377
transform -1 0 680 0 -1 3410
box -4 -6 84 206
use NAND3X1  _3326_
timestamp 1596033377
transform -1 0 744 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3300_
timestamp 1596033377
transform -1 0 808 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3301_
timestamp 1596033377
transform -1 0 856 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3302_
timestamp 1596033377
transform 1 0 856 0 -1 3410
box -4 -6 68 206
use AND2X2  _3243_
timestamp 1596033377
transform -1 0 984 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3370_
timestamp 1596033377
transform 1 0 984 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3371_
timestamp 1596033377
transform 1 0 1048 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3319_
timestamp 1596033377
transform 1 0 1112 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert217
timestamp 1596033377
transform -1 0 1224 0 -1 3410
box -4 -6 52 206
use AND2X2  _3295_
timestamp 1596033377
transform -1 0 1288 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3318_
timestamp 1596033377
transform 1 0 1288 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert216
timestamp 1596033377
transform 1 0 1352 0 -1 3410
box -4 -6 52 206
use FILL  SFILL14000x32100
timestamp 1596033377
transform -1 0 1416 0 -1 3410
box -4 -6 20 206
use AND2X2  _3269_
timestamp 1596033377
transform -1 0 1528 0 -1 3410
box -4 -6 68 206
use AND2X2  _3191_
timestamp 1596033377
transform 1 0 1528 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3270_
timestamp 1596033377
transform -1 0 1656 0 -1 3410
box -4 -6 68 206
use FILL  SFILL14160x32100
timestamp 1596033377
transform -1 0 1432 0 -1 3410
box -4 -6 20 206
use FILL  SFILL14320x32100
timestamp 1596033377
transform -1 0 1448 0 -1 3410
box -4 -6 20 206
use FILL  SFILL14480x32100
timestamp 1596033377
transform -1 0 1464 0 -1 3410
box -4 -6 20 206
use NAND2X1  _3265_
timestamp 1596033377
transform -1 0 1704 0 -1 3410
box -4 -6 52 206
use NOR2X1  _3275_
timestamp 1596033377
transform 1 0 1704 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3274_
timestamp 1596033377
transform -1 0 1816 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3192_
timestamp 1596033377
transform -1 0 1880 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3353_
timestamp 1596033377
transform 1 0 1880 0 -1 3410
box -4 -6 52 206
use NOR2X1  _3223_
timestamp 1596033377
transform 1 0 1928 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3354_
timestamp 1596033377
transform -1 0 2040 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3222_
timestamp 1596033377
transform -1 0 2104 0 -1 3410
box -4 -6 68 206
use INVX1  _3336_
timestamp 1596033377
transform 1 0 2104 0 -1 3410
box -4 -6 36 206
use OAI22X1  _3338_
timestamp 1596033377
transform 1 0 2136 0 -1 3410
box -4 -6 84 206
use INVX1  _3337_
timestamp 1596033377
transform -1 0 2248 0 -1 3410
box -4 -6 36 206
use NOR2X1  _3342_
timestamp 1596033377
transform 1 0 2248 0 -1 3410
box -4 -6 52 206
use OAI21X1  _3341_
timestamp 1596033377
transform 1 0 2296 0 -1 3410
box -4 -6 68 206
use NAND2X1  _3340_
timestamp 1596033377
transform -1 0 2408 0 -1 3410
box -4 -6 52 206
use NAND3X1  _3276_
timestamp 1596033377
transform 1 0 2408 0 -1 3410
box -4 -6 68 206
use NAND3X1  _3224_
timestamp 1596033377
transform -1 0 2536 0 -1 3410
box -4 -6 68 206
use NOR2X1  _3264_
timestamp 1596033377
transform -1 0 2584 0 -1 3410
box -4 -6 52 206
use OAI22X1  _3260_
timestamp 1596033377
transform 1 0 2584 0 -1 3410
box -4 -6 84 206
use INVX1  _3259_
timestamp 1596033377
transform -1 0 2696 0 -1 3410
box -4 -6 36 206
use NOR3X1  _2399_
timestamp 1596033377
transform 1 0 2696 0 -1 3410
box -4 -6 132 206
use NOR2X1  _2388_
timestamp 1596033377
transform -1 0 2872 0 -1 3410
box -4 -6 52 206
use XOR2X1  _2386_
timestamp 1596033377
transform -1 0 3048 0 -1 3410
box -4 -6 116 206
use FILL  SFILL28720x32100
timestamp 1596033377
transform -1 0 2888 0 -1 3410
box -4 -6 20 206
use FILL  SFILL28880x32100
timestamp 1596033377
transform -1 0 2904 0 -1 3410
box -4 -6 20 206
use FILL  SFILL29040x32100
timestamp 1596033377
transform -1 0 2920 0 -1 3410
box -4 -6 20 206
use FILL  SFILL29200x32100
timestamp 1596033377
transform -1 0 2936 0 -1 3410
box -4 -6 20 206
use INVX1  _3206_
timestamp 1596033377
transform -1 0 3080 0 -1 3410
box -4 -6 36 206
use DFFPOSX1  _4572_
timestamp 1596033377
transform -1 0 3272 0 -1 3410
box -4 -6 196 206
use INVX1  _4508_
timestamp 1596033377
transform -1 0 3304 0 -1 3410
box -4 -6 36 206
use NOR2X1  _4507_
timestamp 1596033377
transform -1 0 3352 0 -1 3410
box -4 -6 52 206
use NAND3X1  _4515_
timestamp 1596033377
transform -1 0 3416 0 -1 3410
box -4 -6 68 206
use NAND3X1  _4516_
timestamp 1596033377
transform -1 0 3480 0 -1 3410
box -4 -6 68 206
use NAND2X1  _2127_
timestamp 1596033377
transform -1 0 3528 0 -1 3410
box -4 -6 52 206
use INVX2  _4505_
timestamp 1596033377
transform -1 0 3560 0 -1 3410
box -4 -6 36 206
use OAI21X1  _2137_
timestamp 1596033377
transform 1 0 3560 0 -1 3410
box -4 -6 68 206
use INVX1  _2135_
timestamp 1596033377
transform -1 0 3656 0 -1 3410
box -4 -6 36 206
use AOI21X1  _4518_
timestamp 1596033377
transform 1 0 3656 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4573_
timestamp 1596033377
transform 1 0 3720 0 -1 3410
box -4 -6 196 206
use AOI22X1  _4517_
timestamp 1596033377
transform -1 0 3992 0 -1 3410
box -4 -6 84 206
use OAI21X1  _4616_
timestamp 1596033377
transform -1 0 4056 0 -1 3410
box -4 -6 68 206
use OAI21X1  _4607_
timestamp 1596033377
transform -1 0 4120 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert178
timestamp 1596033377
transform -1 0 4168 0 -1 3410
box -4 -6 52 206
use NOR3X1  _4561_
timestamp 1596033377
transform 1 0 4168 0 -1 3410
box -4 -6 132 206
use OAI21X1  _4610_
timestamp 1596033377
transform -1 0 4360 0 -1 3410
box -4 -6 68 206
use OAI21X1  _4625_
timestamp 1596033377
transform -1 0 4424 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert182
timestamp 1596033377
transform -1 0 4536 0 -1 3410
box -4 -6 52 206
use NOR2X1  _3830_
timestamp 1596033377
transform -1 0 4584 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4388_
timestamp 1596033377
transform 1 0 4584 0 -1 3410
box -4 -6 196 206
use FILL  SFILL44240x32100
timestamp 1596033377
transform -1 0 4440 0 -1 3410
box -4 -6 20 206
use FILL  SFILL44400x32100
timestamp 1596033377
transform -1 0 4456 0 -1 3410
box -4 -6 20 206
use FILL  SFILL44560x32100
timestamp 1596033377
transform -1 0 4472 0 -1 3410
box -4 -6 20 206
use FILL  SFILL44720x32100
timestamp 1596033377
transform -1 0 4488 0 -1 3410
box -4 -6 20 206
use DFFPOSX1  _4308_
timestamp 1596033377
transform 1 0 4776 0 -1 3410
box -4 -6 196 206
use OAI21X1  _3865_
timestamp 1596033377
transform 1 0 4968 0 -1 3410
box -4 -6 68 206
use NAND2X1  _3864_
timestamp 1596033377
transform -1 0 5080 0 -1 3410
box -4 -6 52 206
use NOR2X1  _4288_
timestamp 1596033377
transform 1 0 5080 0 -1 3410
box -4 -6 52 206
use AOI21X1  _4289_
timestamp 1596033377
transform -1 0 5192 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4420_
timestamp 1596033377
transform 1 0 5192 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  _4309_
timestamp 1596033377
transform 1 0 5384 0 -1 3410
box -4 -6 196 206
use OAI21X1  _3867_
timestamp 1596033377
transform 1 0 5576 0 -1 3410
box -4 -6 68 206
use NAND2X1  _3866_
timestamp 1596033377
transform -1 0 5688 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert221
timestamp 1596033377
transform -1 0 5736 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4419_
timestamp 1596033377
transform 1 0 5736 0 -1 3410
box -4 -6 196 206
use DFFPOSX1  _4403_
timestamp 1596033377
transform -1 0 6184 0 -1 3410
box -4 -6 196 206
use FILL  SFILL59280x32100
timestamp 1596033377
transform -1 0 5944 0 -1 3410
box -4 -6 20 206
use FILL  SFILL59440x32100
timestamp 1596033377
transform -1 0 5960 0 -1 3410
box -4 -6 20 206
use FILL  SFILL59600x32100
timestamp 1596033377
transform -1 0 5976 0 -1 3410
box -4 -6 20 206
use FILL  SFILL59760x32100
timestamp 1596033377
transform -1 0 5992 0 -1 3410
box -4 -6 20 206
use DFFPOSX1  _4336_
timestamp 1596033377
transform -1 0 6376 0 -1 3410
box -4 -6 196 206
use NOR2X1  _3889_
timestamp 1596033377
transform 1 0 6376 0 -1 3410
box -4 -6 52 206
use AOI21X1  _3890_
timestamp 1596033377
transform -1 0 6488 0 -1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert255
timestamp 1596033377
transform 1 0 6488 0 -1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert49
timestamp 1596033377
transform 1 0 6536 0 -1 3410
box -4 -6 52 206
use DFFPOSX1  _4379_
timestamp 1596033377
transform -1 0 6776 0 -1 3410
box -4 -6 196 206
use AOI21X1  _3811_
timestamp 1596033377
transform -1 0 6840 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4378_
timestamp 1596033377
transform -1 0 7032 0 -1 3410
box -4 -6 196 206
use OAI21X1  _3796_
timestamp 1596033377
transform 1 0 7032 0 -1 3410
box -4 -6 68 206
use NAND2X1  _3795_
timestamp 1596033377
transform -1 0 7144 0 -1 3410
box -4 -6 52 206
use AOI21X1  _3833_
timestamp 1596033377
transform 1 0 7144 0 -1 3410
box -4 -6 68 206
use DFFPOSX1  _4355_
timestamp 1596033377
transform -1 0 7400 0 -1 3410
box -4 -6 196 206
use INVX1  _3229_
timestamp 1596033377
transform 1 0 8 0 1 3410
box -4 -6 36 206
use OAI22X1  _3230_
timestamp 1596033377
transform -1 0 120 0 1 3410
box -4 -6 84 206
use INVX1  _3333_
timestamp 1596033377
transform 1 0 120 0 1 3410
box -4 -6 36 206
use OAI22X1  _3334_
timestamp 1596033377
transform -1 0 232 0 1 3410
box -4 -6 84 206
use INVX1  _3228_
timestamp 1596033377
transform 1 0 8 0 -1 3810
box -4 -6 36 206
use INVX1  _2557_
timestamp 1596033377
transform -1 0 72 0 -1 3810
box -4 -6 36 206
use AOI21X1  _2558_
timestamp 1596033377
transform -1 0 136 0 -1 3810
box -4 -6 68 206
use AND2X2  _2542_
timestamp 1596033377
transform 1 0 136 0 -1 3810
box -4 -6 68 206
use INVX1  _3332_
timestamp 1596033377
transform -1 0 232 0 -1 3810
box -4 -6 36 206
use INVX1  _3307_
timestamp 1596033377
transform 1 0 232 0 1 3410
box -4 -6 36 206
use OAI22X1  _3308_
timestamp 1596033377
transform -1 0 344 0 1 3410
box -4 -6 84 206
use INVX1  _3306_
timestamp 1596033377
transform -1 0 376 0 1 3410
box -4 -6 36 206
use AND2X2  _2322_
timestamp 1596033377
transform -1 0 440 0 1 3410
box -4 -6 68 206
use NOR2X1  _2550_
timestamp 1596033377
transform -1 0 280 0 -1 3810
box -4 -6 52 206
use XNOR2X1  _2549_
timestamp 1596033377
transform -1 0 392 0 -1 3810
box -4 -6 116 206
use NAND2X1  _2548_
timestamp 1596033377
transform -1 0 440 0 -1 3810
box -4 -6 52 206
use AND2X2  _2365_
timestamp 1596033377
transform 1 0 440 0 1 3410
box -4 -6 68 206
use NAND2X1  _3239_
timestamp 1596033377
transform -1 0 552 0 1 3410
box -4 -6 52 206
use OR2X2  _2354_
timestamp 1596033377
transform 1 0 552 0 1 3410
box -4 -6 68 206
use INVX1  _2546_
timestamp 1596033377
transform -1 0 472 0 -1 3810
box -4 -6 36 206
use INVX1  _3280_
timestamp 1596033377
transform 1 0 472 0 -1 3810
box -4 -6 36 206
use INVX1  _3281_
timestamp 1596033377
transform 1 0 504 0 -1 3810
box -4 -6 36 206
use OAI22X1  _3282_
timestamp 1596033377
transform -1 0 616 0 -1 3810
box -4 -6 84 206
use NOR2X1  _3283_
timestamp 1596033377
transform 1 0 616 0 1 3410
box -4 -6 52 206
use INVX1  _3303_
timestamp 1596033377
transform -1 0 696 0 1 3410
box -4 -6 36 206
use NAND2X1  _3323_
timestamp 1596033377
transform -1 0 744 0 1 3410
box -4 -6 52 206
use AND2X2  _2370_
timestamp 1596033377
transform 1 0 744 0 1 3410
box -4 -6 68 206
use NAND2X1  _3297_
timestamp 1596033377
transform -1 0 856 0 1 3410
box -4 -6 52 206
use INVX1  _3278_
timestamp 1596033377
transform 1 0 616 0 -1 3810
box -4 -6 36 206
use OAI22X1  _3279_
timestamp 1596033377
transform -1 0 728 0 -1 3810
box -4 -6 84 206
use OR2X2  _2352_
timestamp 1596033377
transform -1 0 792 0 -1 3810
box -4 -6 68 206
use AND2X2  _2368_
timestamp 1596033377
transform -1 0 856 0 -1 3810
box -4 -6 68 206
use NOR2X1  _2336_
timestamp 1596033377
transform 1 0 856 0 1 3410
box -4 -6 52 206
use AND2X2  _2337_
timestamp 1596033377
transform 1 0 904 0 1 3410
box -4 -6 68 206
use NOR2X1  _2338_
timestamp 1596033377
transform 1 0 968 0 1 3410
box -4 -6 52 206
use OAI22X1  _3256_
timestamp 1596033377
transform 1 0 856 0 -1 3810
box -4 -6 84 206
use INVX1  _3255_
timestamp 1596033377
transform -1 0 968 0 -1 3810
box -4 -6 36 206
use XOR2X1  _2261_
timestamp 1596033377
transform 1 0 968 0 -1 3810
box -4 -6 116 206
use OAI21X1  _2280_
timestamp 1596033377
transform -1 0 1080 0 1 3410
box -4 -6 68 206
use NAND3X1  _3241_
timestamp 1596033377
transform 1 0 1080 0 1 3410
box -4 -6 68 206
use NAND2X1  _3291_
timestamp 1596033377
transform 1 0 1144 0 1 3410
box -4 -6 52 206
use NAND3X1  _3296_
timestamp 1596033377
transform 1 0 1192 0 1 3410
box -4 -6 68 206
use XNOR2X1  _2262_
timestamp 1596033377
transform -1 0 1192 0 -1 3810
box -4 -6 116 206
use NAND3X1  _3293_
timestamp 1596033377
transform -1 0 1256 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert270
timestamp 1596033377
transform 1 0 1256 0 1 3410
box -4 -6 52 206
use NAND3X1  _3292_
timestamp 1596033377
transform -1 0 1368 0 1 3410
box -4 -6 68 206
use NAND3X1  _3215_
timestamp 1596033377
transform 1 0 1368 0 1 3410
box -4 -6 68 206
use NAND3X1  _3267_
timestamp 1596033377
transform 1 0 1256 0 -1 3810
box -4 -6 68 206
use INVX1  _3176_
timestamp 1596033377
transform 1 0 1320 0 -1 3810
box -4 -6 36 206
use NAND3X1  _3214_
timestamp 1596033377
transform 1 0 1352 0 -1 3810
box -4 -6 68 206
use FILL  SFILL14640x36100
timestamp 1596033377
transform -1 0 1480 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14480x36100
timestamp 1596033377
transform -1 0 1464 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14320x36100
timestamp 1596033377
transform -1 0 1448 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14160x36100
timestamp 1596033377
transform -1 0 1432 0 -1 3810
box -4 -6 20 206
use FILL  SFILL14800x34100
timestamp 1596033377
transform 1 0 1480 0 1 3410
box -4 -6 20 206
use FILL  SFILL14640x34100
timestamp 1596033377
transform 1 0 1464 0 1 3410
box -4 -6 20 206
use FILL  SFILL14480x34100
timestamp 1596033377
transform 1 0 1448 0 1 3410
box -4 -6 20 206
use FILL  SFILL14320x34100
timestamp 1596033377
transform 1 0 1432 0 1 3410
box -4 -6 20 206
use NAND3X1  _3189_
timestamp 1596033377
transform -1 0 1544 0 -1 3810
box -4 -6 68 206
use NAND3X1  _3345_
timestamp 1596033377
transform -1 0 1608 0 -1 3810
box -4 -6 68 206
use AND2X2  _3217_
timestamp 1596033377
transform 1 0 1496 0 1 3410
box -4 -6 68 206
use NAND3X1  _3266_
timestamp 1596033377
transform -1 0 1672 0 -1 3810
box -4 -6 68 206
use NAND3X1  _3218_
timestamp 1596033377
transform -1 0 1624 0 1 3410
box -4 -6 68 206
use NAND2X1  _3213_
timestamp 1596033377
transform -1 0 1672 0 1 3410
box -4 -6 52 206
use NAND2X1  _3271_
timestamp 1596033377
transform 1 0 1672 0 1 3410
box -4 -6 52 206
use AND2X2  _3347_
timestamp 1596033377
transform 1 0 1720 0 1 3410
box -4 -6 68 206
use NAND3X1  _3348_
timestamp 1596033377
transform -1 0 1848 0 1 3410
box -4 -6 68 206
use OAI22X1  _3204_
timestamp 1596033377
transform 1 0 1672 0 -1 3810
box -4 -6 84 206
use INVX1  _3203_
timestamp 1596033377
transform -1 0 1784 0 -1 3810
box -4 -6 36 206
use NAND3X1  _3344_
timestamp 1596033377
transform -1 0 1848 0 -1 3810
box -4 -6 68 206
use NAND2X1  _3343_
timestamp 1596033377
transform 1 0 1848 0 1 3410
box -4 -6 52 206
use OAI22X1  _3178_
timestamp 1596033377
transform 1 0 1896 0 1 3410
box -4 -6 84 206
use INVX1  _3177_
timestamp 1596033377
transform -1 0 2008 0 1 3410
box -4 -6 36 206
use NOR2X1  _3335_
timestamp 1596033377
transform 1 0 2008 0 1 3410
box -4 -6 52 206
use NAND3X1  _3188_
timestamp 1596033377
transform -1 0 1912 0 -1 3810
box -4 -6 68 206
use NOR2X1  _2333_
timestamp 1596033377
transform -1 0 1960 0 -1 3810
box -4 -6 52 206
use NOR2X1  _2335_
timestamp 1596033377
transform 1 0 1960 0 -1 3810
box -4 -6 52 206
use OR2X2  _2353_
timestamp 1596033377
transform 1 0 2008 0 -1 3810
box -4 -6 68 206
use OAI22X1  _3331_
timestamp 1596033377
transform 1 0 2056 0 1 3410
box -4 -6 84 206
use INVX1  _3330_
timestamp 1596033377
transform -1 0 2168 0 1 3410
box -4 -6 36 206
use NAND2X1  _3349_
timestamp 1596033377
transform -1 0 2216 0 1 3410
box -4 -6 52 206
use INVX1  _3329_
timestamp 1596033377
transform 1 0 2072 0 -1 3810
box -4 -6 36 206
use NOR2X1  _3257_
timestamp 1596033377
transform 1 0 2104 0 -1 3810
box -4 -6 52 206
use INVX1  _3252_
timestamp 1596033377
transform -1 0 2184 0 -1 3810
box -4 -6 36 206
use OAI22X1  _3253_
timestamp 1596033377
transform -1 0 2264 0 -1 3810
box -4 -6 84 206
use NOR2X1  _3179_
timestamp 1596033377
transform 1 0 2216 0 1 3410
box -4 -6 52 206
use INVX1  _3339_
timestamp 1596033377
transform 1 0 2264 0 1 3410
box -4 -6 36 206
use NAND2X1  _3193_
timestamp 1596033377
transform -1 0 2344 0 1 3410
box -4 -6 52 206
use OAI22X1  _3175_
timestamp 1596033377
transform 1 0 2344 0 1 3410
box -4 -6 84 206
use NOR2X1  _3205_
timestamp 1596033377
transform 1 0 2264 0 -1 3810
box -4 -6 52 206
use OAI22X1  _3201_
timestamp 1596033377
transform 1 0 2312 0 -1 3810
box -4 -6 84 206
use INVX1  _3200_
timestamp 1596033377
transform -1 0 2424 0 -1 3810
box -4 -6 36 206
use INVX1  _3174_
timestamp 1596033377
transform -1 0 2456 0 1 3410
box -4 -6 36 206
use NAND2X1  _3219_
timestamp 1596033377
transform -1 0 2504 0 1 3410
box -4 -6 52 206
use INVX1  _3173_
timestamp 1596033377
transform -1 0 2536 0 1 3410
box -4 -6 36 206
use OR2X2  _2347_
timestamp 1596033377
transform -1 0 2600 0 1 3410
box -4 -6 68 206
use INVX1  _3258_
timestamp 1596033377
transform -1 0 2632 0 1 3410
box -4 -6 36 206
use INVX1  _3251_
timestamp 1596033377
transform -1 0 2456 0 -1 3810
box -4 -6 36 206
use XNOR2X1  _2420_
timestamp 1596033377
transform -1 0 2568 0 -1 3810
box -4 -6 116 206
use NAND2X1  _2422_
timestamp 1596033377
transform -1 0 2616 0 -1 3810
box -4 -6 52 206
use XOR2X1  _2398_
timestamp 1596033377
transform 1 0 2632 0 1 3410
box -4 -6 116 206
use XOR2X1  _2387_
timestamp 1596033377
transform 1 0 2744 0 1 3410
box -4 -6 116 206
use XOR2X1  _2397_
timestamp 1596033377
transform -1 0 2728 0 -1 3810
box -4 -6 116 206
use AOI22X1  _2427_
timestamp 1596033377
transform -1 0 2808 0 -1 3810
box -4 -6 84 206
use OR2X2  _2426_
timestamp 1596033377
transform -1 0 2872 0 -1 3810
box -4 -6 68 206
use OR2X2  _2350_
timestamp 1596033377
transform -1 0 2936 0 -1 3810
box -4 -6 68 206
use FILL  SFILL29840x36100
timestamp 1596033377
transform -1 0 3000 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29680x36100
timestamp 1596033377
transform -1 0 2984 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29520x36100
timestamp 1596033377
transform -1 0 2968 0 -1 3810
box -4 -6 20 206
use FILL  SFILL29360x36100
timestamp 1596033377
transform -1 0 2952 0 -1 3810
box -4 -6 20 206
use FILL  SFILL30000x34100
timestamp 1596033377
transform 1 0 3000 0 1 3410
box -4 -6 20 206
use FILL  SFILL29840x34100
timestamp 1596033377
transform 1 0 2984 0 1 3410
box -4 -6 20 206
use FILL  SFILL29680x34100
timestamp 1596033377
transform 1 0 2968 0 1 3410
box -4 -6 20 206
use NOR2X1  _2324_
timestamp 1596033377
transform 1 0 3000 0 -1 3810
box -4 -6 52 206
use XNOR2X1  _2409_
timestamp 1596033377
transform 1 0 2856 0 1 3410
box -4 -6 116 206
use AND2X2  _4521_
timestamp 1596033377
transform -1 0 3096 0 1 3410
box -4 -6 68 206
use OAI21X1  _4520_
timestamp 1596033377
transform -1 0 3160 0 1 3410
box -4 -6 68 206
use NOR3X1  _4525_
timestamp 1596033377
transform -1 0 3288 0 1 3410
box -4 -6 132 206
use NOR2X1  _2326_
timestamp 1596033377
transform 1 0 3048 0 -1 3810
box -4 -6 52 206
use DFFPOSX1  _4574_
timestamp 1596033377
transform -1 0 3288 0 -1 3810
box -4 -6 196 206
use FILL  SFILL30160x34100
timestamp 1596033377
transform 1 0 3016 0 1 3410
box -4 -6 20 206
use OAI21X1  _4513_
timestamp 1596033377
transform 1 0 3288 0 1 3410
box -4 -6 68 206
use INVX1  _4512_
timestamp 1596033377
transform -1 0 3384 0 1 3410
box -4 -6 36 206
use INVX1  _2138_
timestamp 1596033377
transform -1 0 3416 0 1 3410
box -4 -6 36 206
use OAI21X1  _2128_
timestamp 1596033377
transform -1 0 3480 0 1 3410
box -4 -6 68 206
use OAI21X1  _4522_
timestamp 1596033377
transform 1 0 3288 0 -1 3810
box -4 -6 68 206
use AOI21X1  _4524_
timestamp 1596033377
transform -1 0 3416 0 -1 3810
box -4 -6 68 206
use NAND3X1  _4526_
timestamp 1596033377
transform -1 0 3480 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4576_
timestamp 1596033377
transform -1 0 3672 0 1 3410
box -4 -6 196 206
use AOI22X1  _4523_
timestamp 1596033377
transform -1 0 3560 0 -1 3810
box -4 -6 84 206
use NAND3X1  _4529_
timestamp 1596033377
transform -1 0 3624 0 -1 3810
box -4 -6 68 206
use AND2X2  _4538_
timestamp 1596033377
transform -1 0 3736 0 1 3410
box -4 -6 68 206
use OAI21X1  _4535_
timestamp 1596033377
transform 1 0 3736 0 1 3410
box -4 -6 68 206
use OAI21X1  _4537_
timestamp 1596033377
transform 1 0 3800 0 1 3410
box -4 -6 68 206
use AOI21X1  _4531_
timestamp 1596033377
transform 1 0 3624 0 -1 3810
box -4 -6 68 206
use AOI22X1  _4530_
timestamp 1596033377
transform -1 0 3768 0 -1 3810
box -4 -6 84 206
use NOR2X1  _4533_
timestamp 1596033377
transform -1 0 3816 0 -1 3810
box -4 -6 52 206
use INVX1  _4532_
timestamp 1596033377
transform -1 0 3848 0 -1 3810
box -4 -6 36 206
use NAND2X1  _4615_
timestamp 1596033377
transform -1 0 3912 0 1 3410
box -4 -6 52 206
use AOI22X1  _4536_
timestamp 1596033377
transform -1 0 3992 0 1 3410
box -4 -6 84 206
use NAND2X1  _4609_
timestamp 1596033377
transform -1 0 4040 0 1 3410
box -4 -6 52 206
use OAI21X1  _4613_
timestamp 1596033377
transform -1 0 3912 0 -1 3810
box -4 -6 68 206
use NAND3X1  _4546_
timestamp 1596033377
transform 1 0 3912 0 -1 3810
box -4 -6 68 206
use AOI22X1  _4542_
timestamp 1596033377
transform -1 0 4056 0 -1 3810
box -4 -6 84 206
use NAND2X1  _4606_
timestamp 1596033377
transform 1 0 4040 0 1 3410
box -4 -6 52 206
use NAND3X1  _4555_
timestamp 1596033377
transform 1 0 4088 0 1 3410
box -4 -6 68 206
use OAI21X1  _4554_
timestamp 1596033377
transform 1 0 4152 0 1 3410
box -4 -6 68 206
use NAND2X1  _4624_
timestamp 1596033377
transform -1 0 4264 0 1 3410
box -4 -6 52 206
use NAND3X1  _4552_
timestamp 1596033377
transform -1 0 4120 0 -1 3810
box -4 -6 68 206
use NOR2X1  _4547_
timestamp 1596033377
transform -1 0 4168 0 -1 3810
box -4 -6 52 206
use INVX1  _4545_
timestamp 1596033377
transform 1 0 4168 0 -1 3810
box -4 -6 36 206
use INVX1  _4553_
timestamp 1596033377
transform -1 0 4232 0 -1 3810
box -4 -6 36 206
use CLKBUF1  CLKBUF1_insert23
timestamp 1596033377
transform -1 0 4408 0 1 3410
box -4 -6 148 206
use AOI22X1  _4549_
timestamp 1596033377
transform -1 0 4312 0 -1 3810
box -4 -6 84 206
use AOI22X1  _4556_
timestamp 1596033377
transform -1 0 4392 0 -1 3810
box -4 -6 84 206
use AOI21X1  _4557_
timestamp 1596033377
transform 1 0 4392 0 -1 3810
box -4 -6 68 206
use FILL  SFILL44080x34100
timestamp 1596033377
transform 1 0 4408 0 1 3410
box -4 -6 20 206
use FILL  SFILL45040x36100
timestamp 1596033377
transform -1 0 4520 0 -1 3810
box -4 -6 20 206
use FILL  SFILL44880x36100
timestamp 1596033377
transform -1 0 4504 0 -1 3810
box -4 -6 20 206
use FILL  SFILL44720x36100
timestamp 1596033377
transform -1 0 4488 0 -1 3810
box -4 -6 20 206
use FILL  SFILL44560x36100
timestamp 1596033377
transform -1 0 4472 0 -1 3810
box -4 -6 20 206
use FILL  SFILL44560x34100
timestamp 1596033377
transform 1 0 4456 0 1 3410
box -4 -6 20 206
use FILL  SFILL44400x34100
timestamp 1596033377
transform 1 0 4440 0 1 3410
box -4 -6 20 206
use FILL  SFILL44240x34100
timestamp 1596033377
transform 1 0 4424 0 1 3410
box -4 -6 20 206
use AOI21X1  _3831_
timestamp 1596033377
transform 1 0 4472 0 1 3410
box -4 -6 68 206
use OAI21X1  _4622_
timestamp 1596033377
transform -1 0 4648 0 -1 3810
box -4 -6 68 206
use OAI21X1  _4619_
timestamp 1596033377
transform -1 0 4584 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4356_
timestamp 1596033377
transform -1 0 4728 0 1 3410
box -4 -6 196 206
use NAND2X1  _3797_
timestamp 1596033377
transform 1 0 4728 0 1 3410
box -4 -6 52 206
use OAI21X1  _3798_
timestamp 1596033377
transform -1 0 4840 0 1 3410
box -4 -6 68 206
use AOI21X1  _3898_
timestamp 1596033377
transform 1 0 4648 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4372_
timestamp 1596033377
transform 1 0 4712 0 -1 3810
box -4 -6 196 206
use MUX2X1  _4219_
timestamp 1596033377
transform 1 0 4840 0 1 3410
box -4 -6 100 206
use MUX2X1  _4041_
timestamp 1596033377
transform -1 0 5032 0 1 3410
box -4 -6 100 206
use OAI21X1  _3731_
timestamp 1596033377
transform 1 0 4904 0 -1 3810
box -4 -6 68 206
use OAI21X1  _3730_
timestamp 1596033377
transform -1 0 5032 0 -1 3810
box -4 -6 68 206
use MUX2X1  _4223_
timestamp 1596033377
transform -1 0 5128 0 1 3410
box -4 -6 100 206
use DFFPOSX1  _4404_
timestamp 1596033377
transform -1 0 5320 0 1 3410
box -4 -6 196 206
use OAI22X1  _4226_
timestamp 1596033377
transform -1 0 5112 0 -1 3810
box -4 -6 84 206
use NOR2X1  _4224_
timestamp 1596033377
transform 1 0 5112 0 -1 3810
box -4 -6 52 206
use OAI21X1  _4225_
timestamp 1596033377
transform -1 0 5224 0 -1 3810
box -4 -6 68 206
use MUX2X1  _4045_
timestamp 1596033377
transform -1 0 5416 0 1 3410
box -4 -6 100 206
use AOI21X1  _3689_
timestamp 1596033377
transform 1 0 5416 0 1 3410
box -4 -6 68 206
use OAI21X1  _4047_
timestamp 1596033377
transform 1 0 5224 0 -1 3810
box -4 -6 68 206
use NOR2X1  _4046_
timestamp 1596033377
transform 1 0 5288 0 -1 3810
box -4 -6 52 206
use OAI22X1  _4048_
timestamp 1596033377
transform 1 0 5336 0 -1 3810
box -4 -6 84 206
use OAI21X1  _4043_
timestamp 1596033377
transform -1 0 5480 0 -1 3810
box -4 -6 68 206
use NOR2X1  _3688_
timestamp 1596033377
transform 1 0 5480 0 1 3410
box -4 -6 52 206
use NOR2X1  _4286_
timestamp 1596033377
transform -1 0 5576 0 1 3410
box -4 -6 52 206
use AOI21X1  _4287_
timestamp 1596033377
transform -1 0 5640 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert67
timestamp 1596033377
transform -1 0 5528 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3869_
timestamp 1596033377
transform -1 0 5592 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert146
timestamp 1596033377
transform -1 0 5640 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert92
timestamp 1596033377
transform -1 0 5688 0 1 3410
box -4 -6 52 206
use AOI21X1  _3686_
timestamp 1596033377
transform 1 0 5688 0 1 3410
box -4 -6 68 206
use NOR2X1  _3685_
timestamp 1596033377
transform -1 0 5800 0 1 3410
box -4 -6 52 206
use MUX2X1  _4034_
timestamp 1596033377
transform 1 0 5800 0 1 3410
box -4 -6 100 206
use NAND2X1  _3763_
timestamp 1596033377
transform 1 0 5640 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3764_
timestamp 1596033377
transform 1 0 5688 0 -1 3810
box -4 -6 68 206
use DFFPOSX1  _4324_
timestamp 1596033377
transform -1 0 5944 0 -1 3810
box -4 -6 196 206
use FILL  SFILL59120x34100
timestamp 1596033377
transform 1 0 5912 0 1 3410
box -4 -6 20 206
use FILL  SFILL58960x34100
timestamp 1596033377
transform 1 0 5896 0 1 3410
box -4 -6 20 206
use FILL  SFILL59920x36100
timestamp 1596033377
transform -1 0 6008 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59760x36100
timestamp 1596033377
transform -1 0 5992 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59600x36100
timestamp 1596033377
transform -1 0 5976 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59440x36100
timestamp 1596033377
transform -1 0 5960 0 -1 3810
box -4 -6 20 206
use FILL  SFILL59440x34100
timestamp 1596033377
transform 1 0 5944 0 1 3410
box -4 -6 20 206
use FILL  SFILL59280x34100
timestamp 1596033377
transform 1 0 5928 0 1 3410
box -4 -6 20 206
use OAI21X1  _4036_
timestamp 1596033377
transform -1 0 6072 0 -1 3810
box -4 -6 68 206
use MUX2X1  _4212_
timestamp 1596033377
transform -1 0 6056 0 1 3410
box -4 -6 100 206
use NOR2X1  _3895_
timestamp 1596033377
transform -1 0 6104 0 1 3410
box -4 -6 52 206
use AOI21X1  _3896_
timestamp 1596033377
transform -1 0 6168 0 1 3410
box -4 -6 68 206
use DFFPOSX1  _4339_
timestamp 1596033377
transform 1 0 6168 0 1 3410
box -4 -6 196 206
use BUFX2  BUFX2_insert13
timestamp 1596033377
transform 1 0 6072 0 -1 3810
box -4 -6 52 206
use OAI21X1  _3863_
timestamp 1596033377
transform -1 0 6184 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert70
timestamp 1596033377
transform 1 0 6184 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert36
timestamp 1596033377
transform -1 0 6408 0 1 3410
box -4 -6 52 206
use DFFPOSX1  _4323_
timestamp 1596033377
transform -1 0 6600 0 1 3410
box -4 -6 196 206
use DFFPOSX1  _4307_
timestamp 1596033377
transform 1 0 6232 0 -1 3810
box -4 -6 196 206
use NAND2X1  _3761_
timestamp 1596033377
transform 1 0 6600 0 1 3410
box -4 -6 52 206
use BUFX2  BUFX2_insert145
timestamp 1596033377
transform 1 0 6424 0 -1 3810
box -4 -6 52 206
use OAI22X1  _4215_
timestamp 1596033377
transform -1 0 6552 0 -1 3810
box -4 -6 84 206
use NOR2X1  _4213_
timestamp 1596033377
transform 1 0 6552 0 -1 3810
box -4 -6 52 206
use OAI21X1  _4214_
timestamp 1596033377
transform 1 0 6600 0 -1 3810
box -4 -6 68 206
use OAI21X1  _3762_
timestamp 1596033377
transform -1 0 6712 0 1 3410
box -4 -6 68 206
use BUFX2  BUFX2_insert7
timestamp 1596033377
transform -1 0 6760 0 1 3410
box -4 -6 52 206
use NOR2X1  _3810_
timestamp 1596033377
transform 1 0 6760 0 1 3410
box -4 -6 52 206
use NOR2X1  _3828_
timestamp 1596033377
transform -1 0 6856 0 1 3410
box -4 -6 52 206
use NOR2X1  _4209_
timestamp 1596033377
transform -1 0 6712 0 -1 3810
box -4 -6 52 206
use OAI21X1  _4210_
timestamp 1596033377
transform 1 0 6712 0 -1 3810
box -4 -6 68 206
use OAI22X1  _4211_
timestamp 1596033377
transform 1 0 6776 0 -1 3810
box -4 -6 84 206
use AOI21X1  _3829_
timestamp 1596033377
transform -1 0 6920 0 1 3410
box -4 -6 68 206
use DFFPOSX1  _4387_
timestamp 1596033377
transform -1 0 7112 0 1 3410
box -4 -6 196 206
use MUX2X1  _4030_
timestamp 1596033377
transform 1 0 6856 0 -1 3810
box -4 -6 100 206
use MUX2X1  _4208_
timestamp 1596033377
transform 1 0 6952 0 -1 3810
box -4 -6 100 206
use AOI21X1  _3823_
timestamp 1596033377
transform 1 0 7112 0 1 3410
box -4 -6 68 206
use DFFPOSX1  _4384_
timestamp 1596033377
transform -1 0 7368 0 1 3410
box -4 -6 196 206
use OAI21X1  _3728_
timestamp 1596033377
transform 1 0 7048 0 -1 3810
box -4 -6 68 206
use OAI21X1  _3729_
timestamp 1596033377
transform 1 0 7112 0 -1 3810
box -4 -6 68 206
use OAI21X1  _3802_
timestamp 1596033377
transform 1 0 7176 0 -1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert51
timestamp 1596033377
transform -1 0 7288 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert50
timestamp 1596033377
transform -1 0 7336 0 -1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert53
timestamp 1596033377
transform -1 0 7384 0 -1 3810
box -4 -6 52 206
use FILL  FILL71120x34100
timestamp 1596033377
transform 1 0 7368 0 1 3410
box -4 -6 20 206
use FILL  FILL71280x34100
timestamp 1596033377
transform 1 0 7384 0 1 3410
box -4 -6 20 206
use FILL  FILL71280x36100
timestamp 1596033377
transform -1 0 7400 0 -1 3810
box -4 -6 20 206
use NAND2X1  _2566_
timestamp 1596033377
transform 1 0 8 0 1 3810
box -4 -6 52 206
use OAI21X1  _2559_
timestamp 1596033377
transform -1 0 120 0 1 3810
box -4 -6 68 206
use XNOR2X1  _2554_
timestamp 1596033377
transform -1 0 232 0 1 3810
box -4 -6 116 206
use AOI21X1  _2552_
timestamp 1596033377
transform -1 0 296 0 1 3810
box -4 -6 68 206
use OAI21X1  _2543_
timestamp 1596033377
transform 1 0 296 0 1 3810
box -4 -6 68 206
use XNOR2X1  _2534_
timestamp 1596033377
transform 1 0 360 0 1 3810
box -4 -6 116 206
use OAI21X1  _2551_
timestamp 1596033377
transform -1 0 536 0 1 3810
box -4 -6 68 206
use NAND2X1  _2533_
timestamp 1596033377
transform -1 0 584 0 1 3810
box -4 -6 52 206
use OR2X2  _2532_
timestamp 1596033377
transform -1 0 648 0 1 3810
box -4 -6 68 206
use NAND2X1  _2531_
timestamp 1596033377
transform -1 0 696 0 1 3810
box -4 -6 52 206
use INVX1  _2530_
timestamp 1596033377
transform -1 0 728 0 1 3810
box -4 -6 36 206
use NOR2X1  _2545_
timestamp 1596033377
transform 1 0 728 0 1 3810
box -4 -6 52 206
use NAND2X1  _2547_
timestamp 1596033377
transform -1 0 824 0 1 3810
box -4 -6 52 206
use INVX1  _2544_
timestamp 1596033377
transform -1 0 856 0 1 3810
box -4 -6 36 206
use AND2X2  _2367_
timestamp 1596033377
transform 1 0 856 0 1 3810
box -4 -6 68 206
use XNOR2X1  _2498_
timestamp 1596033377
transform -1 0 1032 0 1 3810
box -4 -6 116 206
use NAND2X1  _2289_
timestamp 1596033377
transform -1 0 1080 0 1 3810
box -4 -6 52 206
use NAND2X1  _2263_
timestamp 1596033377
transform -1 0 1128 0 1 3810
box -4 -6 52 206
use NOR2X1  _2257_
timestamp 1596033377
transform 1 0 1128 0 1 3810
box -4 -6 52 206
use NOR2X1  _2258_
timestamp 1596033377
transform 1 0 1176 0 1 3810
box -4 -6 52 206
use AOI21X1  _2260_
timestamp 1596033377
transform -1 0 1288 0 1 3810
box -4 -6 68 206
use XOR2X1  _2259_
timestamp 1596033377
transform -1 0 1400 0 1 3810
box -4 -6 116 206
use FILL  SFILL14000x38100
timestamp 1596033377
transform 1 0 1400 0 1 3810
box -4 -6 20 206
use XNOR2X1  _2220_
timestamp 1596033377
transform -1 0 1576 0 1 3810
box -4 -6 116 206
use XNOR2X1  _2273_
timestamp 1596033377
transform -1 0 1688 0 1 3810
box -4 -6 116 206
use FILL  SFILL14160x38100
timestamp 1596033377
transform 1 0 1416 0 1 3810
box -4 -6 20 206
use FILL  SFILL14320x38100
timestamp 1596033377
transform 1 0 1432 0 1 3810
box -4 -6 20 206
use FILL  SFILL14480x38100
timestamp 1596033377
transform 1 0 1448 0 1 3810
box -4 -6 20 206
use NOR2X1  _2330_
timestamp 1596033377
transform -1 0 1736 0 1 3810
box -4 -6 52 206
use NOR2X1  _2332_
timestamp 1596033377
transform 1 0 1736 0 1 3810
box -4 -6 52 206
use AND2X2  _2331_
timestamp 1596033377
transform -1 0 1848 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert1
timestamp 1596033377
transform -1 0 1896 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert242
timestamp 1596033377
transform -1 0 1944 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert243
timestamp 1596033377
transform -1 0 1992 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert41
timestamp 1596033377
transform 1 0 1992 0 1 3810
box -4 -6 52 206
use AND2X2  _2316_
timestamp 1596033377
transform 1 0 2040 0 1 3810
box -4 -6 68 206
use NOR2X1  _2317_
timestamp 1596033377
transform -1 0 2152 0 1 3810
box -4 -6 52 206
use AND2X2  _2334_
timestamp 1596033377
transform -1 0 2216 0 1 3810
box -4 -6 68 206
use AND2X2  _2369_
timestamp 1596033377
transform 1 0 2216 0 1 3810
box -4 -6 68 206
use NOR2X1  _2315_
timestamp 1596033377
transform -1 0 2328 0 1 3810
box -4 -6 52 206
use AND2X2  _2363_
timestamp 1596033377
transform -1 0 2392 0 1 3810
box -4 -6 68 206
use NAND2X1  _2759_
timestamp 1596033377
transform 1 0 2392 0 1 3810
box -4 -6 52 206
use OAI21X1  _2744_
timestamp 1596033377
transform -1 0 2504 0 1 3810
box -4 -6 68 206
use XNOR2X1  _2421_
timestamp 1596033377
transform -1 0 2616 0 1 3810
box -4 -6 116 206
use BUFX2  BUFX2_insert42
timestamp 1596033377
transform 1 0 2616 0 1 3810
box -4 -6 52 206
use AND2X2  _2364_
timestamp 1596033377
transform -1 0 2728 0 1 3810
box -4 -6 68 206
use NAND2X1  _2425_
timestamp 1596033377
transform -1 0 2776 0 1 3810
box -4 -6 52 206
use INVX1  _3199_
timestamp 1596033377
transform -1 0 2808 0 1 3810
box -4 -6 36 206
use OR2X2  _2348_
timestamp 1596033377
transform -1 0 2872 0 1 3810
box -4 -6 68 206
use NAND2X1  _2423_
timestamp 1596033377
transform -1 0 2920 0 1 3810
box -4 -6 52 206
use OR2X2  _2424_
timestamp 1596033377
transform 1 0 2984 0 1 3810
box -4 -6 68 206
use FILL  SFILL29200x38100
timestamp 1596033377
transform 1 0 2920 0 1 3810
box -4 -6 20 206
use FILL  SFILL29360x38100
timestamp 1596033377
transform 1 0 2936 0 1 3810
box -4 -6 20 206
use FILL  SFILL29520x38100
timestamp 1596033377
transform 1 0 2952 0 1 3810
box -4 -6 20 206
use FILL  SFILL29680x38100
timestamp 1596033377
transform 1 0 2968 0 1 3810
box -4 -6 20 206
use BUFX2  BUFX2_insert245
timestamp 1596033377
transform -1 0 3096 0 1 3810
box -4 -6 52 206
use AND2X2  _2325_
timestamp 1596033377
transform -1 0 3160 0 1 3810
box -4 -6 68 206
use BUFX2  BUFX2_insert0
timestamp 1596033377
transform -1 0 3208 0 1 3810
box -4 -6 52 206
use INVX2  _4519_
timestamp 1596033377
transform 1 0 3208 0 1 3810
box -4 -6 36 206
use NOR3X1  _4534_
timestamp 1596033377
transform -1 0 3368 0 1 3810
box -4 -6 132 206
use OAI21X1  _4528_
timestamp 1596033377
transform 1 0 3368 0 1 3810
box -4 -6 68 206
use INVX1  _4527_
timestamp 1596033377
transform -1 0 3464 0 1 3810
box -4 -6 36 206
use DFFPOSX1  _4575_
timestamp 1596033377
transform -1 0 3656 0 1 3810
box -4 -6 196 206
use NOR3X1  _4540_
timestamp 1596033377
transform -1 0 3784 0 1 3810
box -4 -6 132 206
use INVX1  _4539_
timestamp 1596033377
transform -1 0 3816 0 1 3810
box -4 -6 36 206
use NAND2X1  _4612_
timestamp 1596033377
transform -1 0 3864 0 1 3810
box -4 -6 52 206
use OAI21X1  _4541_
timestamp 1596033377
transform 1 0 3864 0 1 3810
box -4 -6 68 206
use OAI21X1  _4543_
timestamp 1596033377
transform 1 0 3928 0 1 3810
box -4 -6 68 206
use AND2X2  _4551_
timestamp 1596033377
transform -1 0 4056 0 1 3810
box -4 -6 68 206
use OAI21X1  _4548_
timestamp 1596033377
transform 1 0 4056 0 1 3810
box -4 -6 68 206
use OAI21X1  _4550_
timestamp 1596033377
transform 1 0 4120 0 1 3810
box -4 -6 68 206
use NAND2X1  _4618_
timestamp 1596033377
transform -1 0 4232 0 1 3810
box -4 -6 52 206
use NAND2X1  _4621_
timestamp 1596033377
transform 1 0 4232 0 1 3810
box -4 -6 52 206
use DFFPOSX1  _4579_
timestamp 1596033377
transform -1 0 4472 0 1 3810
box -4 -6 196 206
use DFFPOSX1  _4340_
timestamp 1596033377
transform -1 0 4728 0 1 3810
box -4 -6 196 206
use FILL  SFILL44720x38100
timestamp 1596033377
transform 1 0 4472 0 1 3810
box -4 -6 20 206
use FILL  SFILL44880x38100
timestamp 1596033377
transform 1 0 4488 0 1 3810
box -4 -6 20 206
use FILL  SFILL45040x38100
timestamp 1596033377
transform 1 0 4504 0 1 3810
box -4 -6 20 206
use FILL  SFILL45200x38100
timestamp 1596033377
transform 1 0 4520 0 1 3810
box -4 -6 20 206
use NOR2X1  _3897_
timestamp 1596033377
transform -1 0 4776 0 1 3810
box -4 -6 52 206
use MUX2X1  _4227_
timestamp 1596033377
transform -1 0 4872 0 1 3810
box -4 -6 100 206
use MUX2X1  _4049_
timestamp 1596033377
transform -1 0 4968 0 1 3810
box -4 -6 100 206
use OAI22X1  _4222_
timestamp 1596033377
transform -1 0 5048 0 1 3810
box -4 -6 84 206
use NOR2X1  _4220_
timestamp 1596033377
transform -1 0 5096 0 1 3810
box -4 -6 52 206
use OAI22X1  _4044_
timestamp 1596033377
transform -1 0 5176 0 1 3810
box -4 -6 84 206
use NOR2X1  _4042_
timestamp 1596033377
transform 1 0 5176 0 1 3810
box -4 -6 52 206
use OAI21X1  _4221_
timestamp 1596033377
transform -1 0 5288 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4310_
timestamp 1596033377
transform -1 0 5480 0 1 3810
box -4 -6 196 206
use NAND2X1  _3868_
timestamp 1596033377
transform 1 0 5480 0 1 3810
box -4 -6 52 206
use DFFPOSX1  _4304_
timestamp 1596033377
transform -1 0 5720 0 1 3810
box -4 -6 196 206
use NAND2X1  _3856_
timestamp 1596033377
transform 1 0 5720 0 1 3810
box -4 -6 52 206
use OAI21X1  _3857_
timestamp 1596033377
transform -1 0 5832 0 1 3810
box -4 -6 68 206
use OAI22X1  _4037_
timestamp 1596033377
transform -1 0 5912 0 1 3810
box -4 -6 84 206
use NOR2X1  _4035_
timestamp 1596033377
transform -1 0 6024 0 1 3810
box -4 -6 52 206
use FILL  SFILL59120x38100
timestamp 1596033377
transform 1 0 5912 0 1 3810
box -4 -6 20 206
use FILL  SFILL59280x38100
timestamp 1596033377
transform 1 0 5928 0 1 3810
box -4 -6 20 206
use FILL  SFILL59440x38100
timestamp 1596033377
transform 1 0 5944 0 1 3810
box -4 -6 20 206
use FILL  SFILL59600x38100
timestamp 1596033377
transform 1 0 5960 0 1 3810
box -4 -6 20 206
use BUFX2  BUFX2_insert276
timestamp 1596033377
transform 1 0 6024 0 1 3810
box -4 -6 52 206
use NAND2X1  _3862_
timestamp 1596033377
transform 1 0 6072 0 1 3810
box -4 -6 52 206
use MUX2X1  _4038_
timestamp 1596033377
transform -1 0 6216 0 1 3810
box -4 -6 100 206
use BUFX2  BUFX2_insert122
timestamp 1596033377
transform 1 0 6216 0 1 3810
box -4 -6 52 206
use MUX2X1  _4216_
timestamp 1596033377
transform -1 0 6360 0 1 3810
box -4 -6 100 206
use OAI22X1  _4033_
timestamp 1596033377
transform -1 0 6440 0 1 3810
box -4 -6 84 206
use OAI21X1  _4032_
timestamp 1596033377
transform -1 0 6504 0 1 3810
box -4 -6 68 206
use NOR2X1  _4031_
timestamp 1596033377
transform -1 0 6552 0 1 3810
box -4 -6 52 206
use MUX2X1  _4175_
timestamp 1596033377
transform -1 0 6648 0 1 3810
box -4 -6 100 206
use MUX2X1  _3997_
timestamp 1596033377
transform 1 0 6648 0 1 3810
box -4 -6 100 206
use NAND2X1  _3789_
timestamp 1596033377
transform 1 0 6744 0 1 3810
box -4 -6 52 206
use OAI21X1  _3790_
timestamp 1596033377
transform -1 0 6856 0 1 3810
box -4 -6 68 206
use DFFPOSX1  _4352_
timestamp 1596033377
transform -1 0 7048 0 1 3810
box -4 -6 196 206
use NOR2X1  _3834_
timestamp 1596033377
transform 1 0 7048 0 1 3810
box -4 -6 52 206
use BUFX2  BUFX2_insert5
timestamp 1596033377
transform 1 0 7096 0 1 3810
box -4 -6 52 206
use NAND2X1  _3801_
timestamp 1596033377
transform 1 0 7144 0 1 3810
box -4 -6 52 206
use DFFPOSX1  _4358_
timestamp 1596033377
transform -1 0 7384 0 1 3810
box -4 -6 196 206
use FILL  FILL71280x38100
timestamp 1596033377
transform 1 0 7384 0 1 3810
box -4 -6 20 206
use NAND3X1  _2562_
timestamp 1596033377
transform -1 0 72 0 -1 4210
box -4 -6 68 206
use INVX1  _2561_
timestamp 1596033377
transform -1 0 104 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2565_
timestamp 1596033377
transform 1 0 104 0 -1 4210
box -4 -6 52 206
use INVX1  _2563_
timestamp 1596033377
transform 1 0 152 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2564_
timestamp 1596033377
transform 1 0 184 0 -1 4210
box -4 -6 68 206
use OAI21X1  _2529_
timestamp 1596033377
transform -1 0 312 0 -1 4210
box -4 -6 68 206
use OR2X2  _2524_
timestamp 1596033377
transform -1 0 376 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2540_
timestamp 1596033377
transform 1 0 376 0 -1 4210
box -4 -6 52 206
use XOR2X1  _2560_
timestamp 1596033377
transform 1 0 424 0 -1 4210
box -4 -6 116 206
use INVX1  _3277_
timestamp 1596033377
transform -1 0 568 0 -1 4210
box -4 -6 36 206
use OR2X2  _2351_
timestamp 1596033377
transform -1 0 632 0 -1 4210
box -4 -6 68 206
use XNOR2X1  _2283_
timestamp 1596033377
transform 1 0 632 0 -1 4210
box -4 -6 116 206
use BUFX2  BUFX2_insert100
timestamp 1596033377
transform -1 0 792 0 -1 4210
box -4 -6 52 206
use AOI21X1  _2281_
timestamp 1596033377
transform 1 0 792 0 -1 4210
box -4 -6 68 206
use INVX1  _2264_
timestamp 1596033377
transform 1 0 856 0 -1 4210
box -4 -6 36 206
use AOI21X1  _2269_
timestamp 1596033377
transform 1 0 888 0 -1 4210
box -4 -6 68 206
use OAI21X1  _2282_
timestamp 1596033377
transform 1 0 952 0 -1 4210
box -4 -6 68 206
use INVX1  _2284_
timestamp 1596033377
transform 1 0 1016 0 -1 4210
box -4 -6 36 206
use NAND3X1  _2285_
timestamp 1596033377
transform 1 0 1048 0 -1 4210
box -4 -6 68 206
use INVX1  _3202_
timestamp 1596033377
transform 1 0 1112 0 -1 4210
box -4 -6 36 206
use BUFX2  BUFX2_insert45
timestamp 1596033377
transform -1 0 1192 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert108
timestamp 1596033377
transform -1 0 1240 0 -1 4210
box -4 -6 52 206
use INVX1  _2266_
timestamp 1596033377
transform -1 0 1272 0 -1 4210
box -4 -6 36 206
use OAI21X1  _2268_
timestamp 1596033377
transform 1 0 1272 0 -1 4210
box -4 -6 68 206
use INVX1  _2265_
timestamp 1596033377
transform -1 0 1368 0 -1 4210
box -4 -6 36 206
use NOR2X1  _2329_
timestamp 1596033377
transform -1 0 1416 0 -1 4210
box -4 -6 52 206
use INVX1  _2593_
timestamp 1596033377
transform -1 0 1512 0 -1 4210
box -4 -6 36 206
use AOI22X1  _2655_
timestamp 1596033377
transform 1 0 1512 0 -1 4210
box -4 -6 84 206
use XNOR2X1  _2569_
timestamp 1596033377
transform 1 0 1592 0 -1 4210
box -4 -6 116 206
use FILL  SFILL14160x40100
timestamp 1596033377
transform -1 0 1432 0 -1 4210
box -4 -6 20 206
use FILL  SFILL14320x40100
timestamp 1596033377
transform -1 0 1448 0 -1 4210
box -4 -6 20 206
use FILL  SFILL14480x40100
timestamp 1596033377
transform -1 0 1464 0 -1 4210
box -4 -6 20 206
use FILL  SFILL14640x40100
timestamp 1596033377
transform -1 0 1480 0 -1 4210
box -4 -6 20 206
use NAND2X1  _2568_
timestamp 1596033377
transform 1 0 1704 0 -1 4210
box -4 -6 52 206
use OAI21X1  _2650_
timestamp 1596033377
transform -1 0 1816 0 -1 4210
box -4 -6 68 206
use NOR2X1  _2648_
timestamp 1596033377
transform 1 0 1816 0 -1 4210
box -4 -6 52 206
use INVX1  _2567_
timestamp 1596033377
transform -1 0 1896 0 -1 4210
box -4 -6 36 206
use BUFX2  BUFX2_insert101
timestamp 1596033377
transform -1 0 1944 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert48
timestamp 1596033377
transform 1 0 1944 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert175
timestamp 1596033377
transform 1 0 1992 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert60
timestamp 1596033377
transform -1 0 2088 0 -1 4210
box -4 -6 52 206
use INVX1  _2656_
timestamp 1596033377
transform -1 0 2120 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2659_
timestamp 1596033377
transform 1 0 2120 0 -1 4210
box -4 -6 52 206
use INVX1  _2658_
timestamp 1596033377
transform -1 0 2200 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2737_
timestamp 1596033377
transform 1 0 2200 0 -1 4210
box -4 -6 52 206
use INVX1  _2745_
timestamp 1596033377
transform 1 0 2248 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2657_
timestamp 1596033377
transform -1 0 2328 0 -1 4210
box -4 -6 52 206
use AOI22X1  _2758_
timestamp 1596033377
transform 1 0 2328 0 -1 4210
box -4 -6 84 206
use AOI22X1  _2739_
timestamp 1596033377
transform 1 0 2408 0 -1 4210
box -4 -6 84 206
use OAI22X1  _2746_
timestamp 1596033377
transform -1 0 2568 0 -1 4210
box -4 -6 84 206
use NAND2X1  _2738_
timestamp 1596033377
transform 1 0 2568 0 -1 4210
box -4 -6 52 206
use AOI21X1  _2747_
timestamp 1596033377
transform -1 0 2680 0 -1 4210
box -4 -6 68 206
use NAND2X1  _2666_
timestamp 1596033377
transform 1 0 2680 0 -1 4210
box -4 -6 52 206
use OAI22X1  _2665_
timestamp 1596033377
transform 1 0 2728 0 -1 4210
box -4 -6 84 206
use INVX1  _2663_
timestamp 1596033377
transform -1 0 2840 0 -1 4210
box -4 -6 36 206
use INVX1  _2664_
timestamp 1596033377
transform 1 0 2840 0 -1 4210
box -4 -6 36 206
use NAND2X1  _2669_
timestamp 1596033377
transform -1 0 2920 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert246
timestamp 1596033377
transform 1 0 2984 0 -1 4210
box -4 -6 52 206
use FILL  SFILL29200x40100
timestamp 1596033377
transform -1 0 2936 0 -1 4210
box -4 -6 20 206
use FILL  SFILL29360x40100
timestamp 1596033377
transform -1 0 2952 0 -1 4210
box -4 -6 20 206
use FILL  SFILL29520x40100
timestamp 1596033377
transform -1 0 2968 0 -1 4210
box -4 -6 20 206
use FILL  SFILL29680x40100
timestamp 1596033377
transform -1 0 2984 0 -1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert110
timestamp 1596033377
transform -1 0 3080 0 -1 4210
box -4 -6 52 206
use XNOR2X1  _2402_
timestamp 1596033377
transform 1 0 3080 0 -1 4210
box -4 -6 116 206
use NAND2X1  _2404_
timestamp 1596033377
transform 1 0 3192 0 -1 4210
box -4 -6 52 206
use NAND2X1  _2157_
timestamp 1596033377
transform -1 0 3288 0 -1 4210
box -4 -6 52 206
use NAND2X1  _2139_
timestamp 1596033377
transform 1 0 3288 0 -1 4210
box -4 -6 52 206
use OAI21X1  _2140_
timestamp 1596033377
transform -1 0 3400 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert198
timestamp 1596033377
transform -1 0 3448 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4050_
timestamp 1596033377
transform 1 0 3448 0 -1 4210
box -4 -6 68 206
use AOI21X1  _4051_
timestamp 1596033377
transform -1 0 3576 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert137
timestamp 1596033377
transform -1 0 3624 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert62
timestamp 1596033377
transform 1 0 3624 0 -1 4210
box -4 -6 52 206
use AOI21X1  _4218_
timestamp 1596033377
transform -1 0 3736 0 -1 4210
box -4 -6 68 206
use NAND2X1  _2151_
timestamp 1596033377
transform -1 0 3784 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert199
timestamp 1596033377
transform -1 0 3832 0 -1 4210
box -4 -6 52 206
use AND2X2  _4544_
timestamp 1596033377
transform -1 0 3896 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4578_
timestamp 1596033377
transform 1 0 3896 0 -1 4210
box -4 -6 196 206
use OAI21X1  _4228_
timestamp 1596033377
transform 1 0 4088 0 -1 4210
box -4 -6 68 206
use AOI21X1  _4229_
timestamp 1596033377
transform -1 0 4216 0 -1 4210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_insert31
timestamp 1596033377
transform -1 0 4360 0 -1 4210
box -4 -6 148 206
use INVX4  _3678_
timestamp 1596033377
transform -1 0 4408 0 -1 4210
box -4 -6 52 206
use FILL  SFILL44080x40100
timestamp 1596033377
transform -1 0 4424 0 -1 4210
box -4 -6 20 206
use AOI21X1  _3825_
timestamp 1596033377
transform 1 0 4472 0 -1 4210
box -4 -6 68 206
use NOR2X1  _3824_
timestamp 1596033377
transform -1 0 4584 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4353_
timestamp 1596033377
transform -1 0 4776 0 -1 4210
box -4 -6 196 206
use FILL  SFILL44240x40100
timestamp 1596033377
transform -1 0 4440 0 -1 4210
box -4 -6 20 206
use FILL  SFILL44400x40100
timestamp 1596033377
transform -1 0 4456 0 -1 4210
box -4 -6 20 206
use FILL  SFILL44560x40100
timestamp 1596033377
transform -1 0 4472 0 -1 4210
box -4 -6 20 206
use NAND2X1  _3791_
timestamp 1596033377
transform 1 0 4776 0 -1 4210
box -4 -6 52 206
use OAI21X1  _3792_
timestamp 1596033377
transform -1 0 4888 0 -1 4210
box -4 -6 68 206
use NOR2X1  _3694_
timestamp 1596033377
transform -1 0 4936 0 -1 4210
box -4 -6 52 206
use AOI21X1  _3695_
timestamp 1596033377
transform -1 0 5000 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4406_
timestamp 1596033377
transform 1 0 5000 0 -1 4210
box -4 -6 196 206
use BUFX2  BUFX2_insert285
timestamp 1596033377
transform -1 0 5240 0 -1 4210
box -4 -6 52 206
use OAI21X1  _4181_
timestamp 1596033377
transform -1 0 5304 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert121
timestamp 1596033377
transform -1 0 5352 0 -1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert275
timestamp 1596033377
transform -1 0 5400 0 -1 4210
box -4 -6 52 206
use DFFPOSX1  _4368_
timestamp 1596033377
transform -1 0 5592 0 -1 4210
box -4 -6 196 206
use OAI21X1  _3723_
timestamp 1596033377
transform 1 0 5592 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3722_
timestamp 1596033377
transform -1 0 5720 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert283
timestamp 1596033377
transform 1 0 5720 0 -1 4210
box -4 -6 52 206
use NOR2X1  _3998_
timestamp 1596033377
transform 1 0 5768 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4000_
timestamp 1596033377
transform 1 0 5816 0 -1 4210
box -4 -6 84 206
use OAI21X1  _3999_
timestamp 1596033377
transform -1 0 5960 0 -1 4210
box -4 -6 68 206
use FILL  SFILL59600x40100
timestamp 1596033377
transform -1 0 5976 0 -1 4210
box -4 -6 20 206
use FILL  SFILL59760x40100
timestamp 1596033377
transform -1 0 5992 0 -1 4210
box -4 -6 20 206
use FILL  SFILL59920x40100
timestamp 1596033377
transform -1 0 6008 0 -1 4210
box -4 -6 20 206
use FILL  SFILL60080x40100
timestamp 1596033377
transform -1 0 6024 0 -1 4210
box -4 -6 20 206
use NOR2X1  _4176_
timestamp 1596033377
transform 1 0 6024 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4178_
timestamp 1596033377
transform 1 0 6072 0 -1 4210
box -4 -6 84 206
use OAI21X1  _4177_
timestamp 1596033377
transform -1 0 6216 0 -1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert210
timestamp 1596033377
transform 1 0 6216 0 -1 4210
box -4 -6 52 206
use NOR2X1  _4242_
timestamp 1596033377
transform -1 0 6312 0 -1 4210
box -4 -6 52 206
use OAI22X1  _4244_
timestamp 1596033377
transform 1 0 6312 0 -1 4210
box -4 -6 84 206
use OAI21X1  _4243_
timestamp 1596033377
transform -1 0 6456 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3734_
timestamp 1596033377
transform 1 0 6456 0 -1 4210
box -4 -6 68 206
use OAI21X1  _3735_
timestamp 1596033377
transform -1 0 6584 0 -1 4210
box -4 -6 68 206
use DFFPOSX1  _4374_
timestamp 1596033377
transform -1 0 6776 0 -1 4210
box -4 -6 196 206
use MUX2X1  _4063_
timestamp 1596033377
transform 1 0 6776 0 -1 4210
box -4 -6 100 206
use MUX2X1  _4241_
timestamp 1596033377
transform -1 0 6968 0 -1 4210
box -4 -6 100 206
use DFFPOSX1  _4326_
timestamp 1596033377
transform -1 0 7160 0 -1 4210
box -4 -6 196 206
use DFFPOSX1  _4390_
timestamp 1596033377
transform -1 0 7352 0 -1 4210
box -4 -6 196 206
use FILL  FILL70960x40100
timestamp 1596033377
transform -1 0 7368 0 -1 4210
box -4 -6 20 206
use FILL  FILL71120x40100
timestamp 1596033377
transform -1 0 7384 0 -1 4210
box -4 -6 20 206
use FILL  FILL71280x40100
timestamp 1596033377
transform -1 0 7400 0 -1 4210
box -4 -6 20 206
use AND2X2  _2514_
timestamp 1596033377
transform -1 0 72 0 1 4210
box -4 -6 68 206
use OR2X2  _2513_
timestamp 1596033377
transform -1 0 136 0 1 4210
box -4 -6 68 206
use NAND2X1  _2512_
timestamp 1596033377
transform -1 0 184 0 1 4210
box -4 -6 52 206
use NAND2X1  _2523_
timestamp 1596033377
transform 1 0 184 0 1 4210
box -4 -6 52 206
use AOI21X1  _2528_
timestamp 1596033377
transform -1 0 296 0 1 4210
box -4 -6 68 206
use INVX1  _2525_
timestamp 1596033377
transform -1 0 328 0 1 4210
box -4 -6 36 206
use INVX1  _2508_
timestamp 1596033377
transform -1 0 360 0 1 4210
box -4 -6 36 206
use OAI21X1  _2510_
timestamp 1596033377
transform -1 0 424 0 1 4210
box -4 -6 68 206
use INVX1  _2555_
timestamp 1596033377
transform 1 0 424 0 1 4210
box -4 -6 36 206
use NAND2X1  _2556_
timestamp 1596033377
transform -1 0 504 0 1 4210
box -4 -6 52 206
use XNOR2X1  _2553_
timestamp 1596033377
transform -1 0 616 0 1 4210
box -4 -6 116 206
use NAND2X1  _2509_
timestamp 1596033377
transform -1 0 664 0 1 4210
box -4 -6 52 206
use OAI21X1  _2500_
timestamp 1596033377
transform -1 0 728 0 1 4210
box -4 -6 68 206
use INVX1  _2499_
timestamp 1596033377
transform -1 0 760 0 1 4210
box -4 -6 36 206
use XOR2X1  _2506_
timestamp 1596033377
transform -1 0 872 0 1 4210
box -4 -6 116 206
use OAI21X1  _2255_
timestamp 1596033377
transform 1 0 872 0 1 4210
box -4 -6 68 206
use AND2X2  _2497_
timestamp 1596033377
transform -1 0 1000 0 1 4210
box -4 -6 68 206
use NAND2X1  _2288_
timestamp 1596033377
transform 1 0 1000 0 1 4210
box -4 -6 52 206
use OAI21X1  _2287_
timestamp 1596033377
transform -1 0 1112 0 1 4210
box -4 -6 68 206
use INVX1  _2286_
timestamp 1596033377
transform -1 0 1144 0 1 4210
box -4 -6 36 206
use NAND2X1  _2270_
timestamp 1596033377
transform -1 0 1192 0 1 4210
box -4 -6 52 206
use AND2X2  _2272_
timestamp 1596033377
transform -1 0 1256 0 1 4210
box -4 -6 68 206
use OR2X2  _2271_
timestamp 1596033377
transform -1 0 1320 0 1 4210
box -4 -6 68 206
use OAI21X1  _2267_
timestamp 1596033377
transform -1 0 1384 0 1 4210
box -4 -6 68 206
use AND2X2  _2328_
timestamp 1596033377
transform -1 0 1448 0 1 4210
box -4 -6 68 206
use OAI21X1  _2653_
timestamp 1596033377
transform 1 0 1512 0 1 4210
box -4 -6 68 206
use NAND2X1  _2654_
timestamp 1596033377
transform -1 0 1624 0 1 4210
box -4 -6 52 206
use FILL  SFILL14480x42100
timestamp 1596033377
transform 1 0 1448 0 1 4210
box -4 -6 20 206
use FILL  SFILL14640x42100
timestamp 1596033377
transform 1 0 1464 0 1 4210
box -4 -6 20 206
use FILL  SFILL14800x42100
timestamp 1596033377
transform 1 0 1480 0 1 4210
box -4 -6 20 206
use FILL  SFILL14960x42100
timestamp 1596033377
transform 1 0 1496 0 1 4210
box -4 -6 20 206
use NOR2X1  _2327_
timestamp 1596033377
transform -1 0 1672 0 1 4210
box -4 -6 52 206
use NAND3X1  _2573_
timestamp 1596033377
transform -1 0 1736 0 1 4210
box -4 -6 68 206
use NAND2X1  _2572_
timestamp 1596033377
transform 1 0 1736 0 1 4210
box -4 -6 52 206
use NOR2X1  _2649_
timestamp 1596033377
transform -1 0 1832 0 1 4210
box -4 -6 52 206
use OR2X2  _2571_
timestamp 1596033377
transform -1 0 1896 0 1 4210
box -4 -6 68 206
use INVX1  _2570_
timestamp 1596033377
transform -1 0 1928 0 1 4210
box -4 -6 36 206
use BUFX2  BUFX2_insert154
timestamp 1596033377
transform -1 0 1976 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert152
timestamp 1596033377
transform 1 0 1976 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert61
timestamp 1596033377
transform -1 0 2072 0 1 4210
box -4 -6 52 206
use NAND2X1  _2938_
timestamp 1596033377
transform -1 0 2120 0 1 4210
box -4 -6 52 206
use NAND3X1  _2937_
timestamp 1596033377
transform -1 0 2184 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert59
timestamp 1596033377
transform 1 0 2184 0 1 4210
box -4 -6 52 206
use OAI21X1  _2930_
timestamp 1596033377
transform 1 0 2232 0 1 4210
box -4 -6 68 206
use NAND3X1  _2662_
timestamp 1596033377
transform 1 0 2296 0 1 4210
box -4 -6 68 206
use NAND2X1  _2661_
timestamp 1596033377
transform 1 0 2360 0 1 4210
box -4 -6 52 206
use AOI21X1  _2743_
timestamp 1596033377
transform 1 0 2408 0 1 4210
box -4 -6 68 206
use NAND2X1  _2687_
timestamp 1596033377
transform 1 0 2472 0 1 4210
box -4 -6 52 206
use OAI21X1  _2742_
timestamp 1596033377
transform -1 0 2584 0 1 4210
box -4 -6 68 206
use NAND3X1  _2748_
timestamp 1596033377
transform 1 0 2584 0 1 4210
box -4 -6 68 206
use INVX1  _2740_
timestamp 1596033377
transform -1 0 2680 0 1 4210
box -4 -6 36 206
use OAI21X1  _2741_
timestamp 1596033377
transform 1 0 2680 0 1 4210
box -4 -6 68 206
use NOR3X1  _2671_
timestamp 1596033377
transform 1 0 2744 0 1 4210
box -4 -6 132 206
use NAND3X1  _2670_
timestamp 1596033377
transform 1 0 2872 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert153
timestamp 1596033377
transform 1 0 3000 0 1 4210
box -4 -6 52 206
use FILL  SFILL29360x42100
timestamp 1596033377
transform 1 0 2936 0 1 4210
box -4 -6 20 206
use FILL  SFILL29520x42100
timestamp 1596033377
transform 1 0 2952 0 1 4210
box -4 -6 20 206
use FILL  SFILL29680x42100
timestamp 1596033377
transform 1 0 2968 0 1 4210
box -4 -6 20 206
use FILL  SFILL29840x42100
timestamp 1596033377
transform 1 0 2984 0 1 4210
box -4 -6 20 206
use BUFX2  BUFX2_insert47
timestamp 1596033377
transform -1 0 3096 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4452_
timestamp 1596033377
transform -1 0 3288 0 1 4210
box -4 -6 196 206
use OAI21X1  _2158_
timestamp 1596033377
transform -1 0 3352 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert197
timestamp 1596033377
transform -1 0 3400 0 1 4210
box -4 -6 52 206
use BUFX2  _2094_
timestamp 1596033377
transform 1 0 3400 0 1 4210
box -4 -6 52 206
use INVX1  _2156_
timestamp 1596033377
transform -1 0 3480 0 1 4210
box -4 -6 36 206
use OAI21X1  _4250_
timestamp 1596033377
transform 1 0 3480 0 1 4210
box -4 -6 68 206
use BUFX2  _2093_
timestamp 1596033377
transform -1 0 3592 0 1 4210
box -4 -6 52 206
use OAI21X1  _4072_
timestamp 1596033377
transform 1 0 3592 0 1 4210
box -4 -6 68 206
use OAI21X1  _4217_
timestamp 1596033377
transform -1 0 3720 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert172
timestamp 1596033377
transform 1 0 3720 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4577_
timestamp 1596033377
transform 1 0 3768 0 1 4210
box -4 -6 196 206
use INVX1  _2153_
timestamp 1596033377
transform -1 0 3992 0 1 4210
box -4 -6 36 206
use INVX1  _2159_
timestamp 1596033377
transform -1 0 4024 0 1 4210
box -4 -6 36 206
use DFFPOSX1  _4436_
timestamp 1596033377
transform -1 0 4216 0 1 4210
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert35
timestamp 1596033377
transform -1 0 4360 0 1 4210
box -4 -6 148 206
use FILL  SFILL43600x42100
timestamp 1596033377
transform 1 0 4360 0 1 4210
box -4 -6 20 206
use FILL  SFILL43760x42100
timestamp 1596033377
transform 1 0 4376 0 1 4210
box -4 -6 20 206
use FILL  SFILL43920x42100
timestamp 1596033377
transform 1 0 4392 0 1 4210
box -4 -6 20 206
use FILL  SFILL44080x42100
timestamp 1596033377
transform 1 0 4408 0 1 4210
box -4 -6 20 206
use DFFPOSX1  _4385_
timestamp 1596033377
transform 1 0 4424 0 1 4210
box -4 -6 196 206
use MUX2X1  _4008_
timestamp 1596033377
transform 1 0 4616 0 1 4210
box -4 -6 100 206
use MUX2X1  _4186_
timestamp 1596033377
transform -1 0 4808 0 1 4210
box -4 -6 100 206
use BUFX2  BUFX2_insert213
timestamp 1596033377
transform 1 0 4808 0 1 4210
box -4 -6 52 206
use INVX4  _3681_
timestamp 1596033377
transform -1 0 4904 0 1 4210
box -4 -6 52 206
use NOR2X1  _4068_
timestamp 1596033377
transform -1 0 4952 0 1 4210
box -4 -6 52 206
use NOR2X1  _4246_
timestamp 1596033377
transform 1 0 4952 0 1 4210
box -4 -6 52 206
use MUX2X1  _4071_
timestamp 1596033377
transform -1 0 5096 0 1 4210
box -4 -6 100 206
use OAI22X1  _4070_
timestamp 1596033377
transform 1 0 5096 0 1 4210
box -4 -6 84 206
use MUX2X1  _4183_
timestamp 1596033377
transform -1 0 5272 0 1 4210
box -4 -6 100 206
use OAI22X1  _4182_
timestamp 1596033377
transform 1 0 5272 0 1 4210
box -4 -6 84 206
use NOR2X1  _4180_
timestamp 1596033377
transform -1 0 5400 0 1 4210
box -4 -6 52 206
use MUX2X1  _4005_
timestamp 1596033377
transform -1 0 5496 0 1 4210
box -4 -6 100 206
use BUFX2  BUFX2_insert259
timestamp 1596033377
transform -1 0 5544 0 1 4210
box -4 -6 52 206
use OAI22X1  _4004_
timestamp 1596033377
transform -1 0 5624 0 1 4210
box -4 -6 84 206
use NOR2X1  _4002_
timestamp 1596033377
transform 1 0 5624 0 1 4210
box -4 -6 52 206
use BUFX2  BUFX2_insert257
timestamp 1596033377
transform -1 0 5720 0 1 4210
box -4 -6 52 206
use OAI21X1  _4003_
timestamp 1596033377
transform 1 0 5720 0 1 4210
box -4 -6 68 206
use OAI21X1  _3732_
timestamp 1596033377
transform 1 0 5784 0 1 4210
box -4 -6 68 206
use OAI21X1  _3733_
timestamp 1596033377
transform -1 0 5912 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4373_
timestamp 1596033377
transform 1 0 5976 0 1 4210
box -4 -6 196 206
use FILL  SFILL59120x42100
timestamp 1596033377
transform 1 0 5912 0 1 4210
box -4 -6 20 206
use FILL  SFILL59280x42100
timestamp 1596033377
transform 1 0 5928 0 1 4210
box -4 -6 20 206
use FILL  SFILL59440x42100
timestamp 1596033377
transform 1 0 5944 0 1 4210
box -4 -6 20 206
use FILL  SFILL59600x42100
timestamp 1596033377
transform 1 0 5960 0 1 4210
box -4 -6 20 206
use NOR2X1  _4064_
timestamp 1596033377
transform -1 0 6216 0 1 4210
box -4 -6 52 206
use OAI22X1  _4066_
timestamp 1596033377
transform 1 0 6216 0 1 4210
box -4 -6 84 206
use OAI21X1  _4065_
timestamp 1596033377
transform -1 0 6360 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4325_
timestamp 1596033377
transform -1 0 6552 0 1 4210
box -4 -6 196 206
use NAND2X1  _3765_
timestamp 1596033377
transform 1 0 6552 0 1 4210
box -4 -6 52 206
use OAI21X1  _3766_
timestamp 1596033377
transform -1 0 6664 0 1 4210
box -4 -6 68 206
use BUFX2  BUFX2_insert40
timestamp 1596033377
transform 1 0 6664 0 1 4210
box -4 -6 52 206
use NAND2X1  _3755_
timestamp 1596033377
transform 1 0 6712 0 1 4210
box -4 -6 52 206
use OAI21X1  _3756_
timestamp 1596033377
transform -1 0 6824 0 1 4210
box -4 -6 68 206
use OAI21X1  _3768_
timestamp 1596033377
transform 1 0 6824 0 1 4210
box -4 -6 68 206
use NAND2X1  _3767_
timestamp 1596033377
transform -1 0 6936 0 1 4210
box -4 -6 52 206
use DFFPOSX1  _4320_
timestamp 1596033377
transform -1 0 7128 0 1 4210
box -4 -6 196 206
use OAI21X1  _3800_
timestamp 1596033377
transform 1 0 7128 0 1 4210
box -4 -6 68 206
use DFFPOSX1  _4357_
timestamp 1596033377
transform -1 0 7384 0 1 4210
box -4 -6 196 206
use FILL  FILL71280x42100
timestamp 1596033377
transform 1 0 7384 0 1 4210
box -4 -6 20 206
use INVX1  _2526_
timestamp 1596033377
transform 1 0 8 0 -1 4610
box -4 -6 36 206
use NOR2X1  _2521_
timestamp 1596033377
transform -1 0 88 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2527_
timestamp 1596033377
transform -1 0 152 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2517_
timestamp 1596033377
transform -1 0 200 0 -1 4610
box -4 -6 52 206
use XOR2X1  _2522_
timestamp 1596033377
transform 1 0 200 0 -1 4610
box -4 -6 116 206
use INVX1  _3254_
timestamp 1596033377
transform 1 0 312 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2247_
timestamp 1596033377
transform 1 0 344 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2246_
timestamp 1596033377
transform 1 0 392 0 -1 4610
box -4 -6 52 206
use INVX1  _2244_
timestamp 1596033377
transform 1 0 440 0 -1 4610
box -4 -6 36 206
use OAI21X1  _2245_
timestamp 1596033377
transform 1 0 472 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2248_
timestamp 1596033377
transform 1 0 536 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2238_
timestamp 1596033377
transform -1 0 632 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2507_
timestamp 1596033377
transform -1 0 696 0 -1 4610
box -4 -6 68 206
use INVX1  _2504_
timestamp 1596033377
transform 1 0 696 0 -1 4610
box -4 -6 36 206
use NOR2X1  _2505_
timestamp 1596033377
transform -1 0 776 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2502_
timestamp 1596033377
transform -1 0 824 0 -1 4610
box -4 -6 52 206
use OR2X2  _2250_
timestamp 1596033377
transform 1 0 824 0 -1 4610
box -4 -6 68 206
use NOR2X1  _2279_
timestamp 1596033377
transform -1 0 936 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2226_
timestamp 1596033377
transform -1 0 984 0 -1 4610
box -4 -6 52 206
use OR2X2  _2496_
timestamp 1596033377
transform -1 0 1048 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2495_
timestamp 1596033377
transform -1 0 1096 0 -1 4610
box -4 -6 52 206
use INVX1  _2494_
timestamp 1596033377
transform -1 0 1128 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2231_
timestamp 1596033377
transform -1 0 1176 0 -1 4610
box -4 -6 52 206
use XOR2X1  _2227_
timestamp 1596033377
transform -1 0 1288 0 -1 4610
box -4 -6 116 206
use BUFX2  BUFX2_insert109
timestamp 1596033377
transform 1 0 1288 0 -1 4610
box -4 -6 52 206
use AND2X2  _2256_
timestamp 1596033377
transform -1 0 1400 0 -1 4610
box -4 -6 68 206
use INVX1  _2645_
timestamp 1596033377
transform 1 0 1400 0 -1 4610
box -4 -6 36 206
use OAI22X1  _2646_
timestamp 1596033377
transform -1 0 1576 0 -1 4610
box -4 -6 84 206
use INVX1  _2644_
timestamp 1596033377
transform -1 0 1608 0 -1 4610
box -4 -6 36 206
use INVX1  _2643_
timestamp 1596033377
transform 1 0 1608 0 -1 4610
box -4 -6 36 206
use FILL  SFILL14320x44100
timestamp 1596033377
transform -1 0 1448 0 -1 4610
box -4 -6 20 206
use FILL  SFILL14480x44100
timestamp 1596033377
transform -1 0 1464 0 -1 4610
box -4 -6 20 206
use FILL  SFILL14640x44100
timestamp 1596033377
transform -1 0 1480 0 -1 4610
box -4 -6 20 206
use FILL  SFILL14800x44100
timestamp 1596033377
transform -1 0 1496 0 -1 4610
box -4 -6 20 206
use OAI21X1  _2647_
timestamp 1596033377
transform 1 0 1640 0 -1 4610
box -4 -6 68 206
use OAI21X1  _2651_
timestamp 1596033377
transform 1 0 1704 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert2
timestamp 1596033377
transform -1 0 1816 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert3
timestamp 1596033377
transform 1 0 1816 0 -1 4610
box -4 -6 52 206
use INVX1  _2856_
timestamp 1596033377
transform 1 0 1864 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2857_
timestamp 1596033377
transform 1 0 1896 0 -1 4610
box -4 -6 52 206
use OAI22X1  _2924_
timestamp 1596033377
transform -1 0 2024 0 -1 4610
box -4 -6 84 206
use INVX1  _2870_
timestamp 1596033377
transform 1 0 2024 0 -1 4610
box -4 -6 36 206
use INVX1  _2858_
timestamp 1596033377
transform 1 0 2056 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2859_
timestamp 1596033377
transform -1 0 2136 0 -1 4610
box -4 -6 52 206
use AND2X2  _2931_
timestamp 1596033377
transform 1 0 2136 0 -1 4610
box -4 -6 68 206
use NAND3X1  _2878_
timestamp 1596033377
transform 1 0 2200 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert195
timestamp 1596033377
transform -1 0 2312 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert46
timestamp 1596033377
transform -1 0 2360 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert192
timestamp 1596033377
transform 1 0 2360 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2750_
timestamp 1596033377
transform 1 0 2408 0 -1 4610
box -4 -6 52 206
use INVX2  _2660_
timestamp 1596033377
transform 1 0 2456 0 -1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert102
timestamp 1596033377
transform 1 0 2488 0 -1 4610
box -4 -6 52 206
use INVX1  _2847_
timestamp 1596033377
transform 1 0 2536 0 -1 4610
box -4 -6 36 206
use AOI21X1  _2927_
timestamp 1596033377
transform 1 0 2568 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2848_
timestamp 1596033377
transform -1 0 2680 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert151
timestamp 1596033377
transform -1 0 2728 0 -1 4610
box -4 -6 52 206
use NOR2X1  _2382_
timestamp 1596033377
transform 1 0 2728 0 -1 4610
box -4 -6 52 206
use OAI22X1  _2383_
timestamp 1596033377
transform -1 0 2856 0 -1 4610
box -4 -6 84 206
use NOR2X1  _2380_
timestamp 1596033377
transform 1 0 2856 0 -1 4610
box -4 -6 52 206
use AND2X2  _2379_
timestamp 1596033377
transform -1 0 3032 0 -1 4610
box -4 -6 68 206
use FILL  SFILL29040x44100
timestamp 1596033377
transform -1 0 2920 0 -1 4610
box -4 -6 20 206
use FILL  SFILL29200x44100
timestamp 1596033377
transform -1 0 2936 0 -1 4610
box -4 -6 20 206
use FILL  SFILL29360x44100
timestamp 1596033377
transform -1 0 2952 0 -1 4610
box -4 -6 20 206
use FILL  SFILL29520x44100
timestamp 1596033377
transform -1 0 2968 0 -1 4610
box -4 -6 20 206
use DFFPOSX1  _4438_
timestamp 1596033377
transform -1 0 3224 0 -1 4610
box -4 -6 196 206
use DFFPOSX1  _4453_
timestamp 1596033377
transform -1 0 3416 0 -1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert194
timestamp 1596033377
transform -1 0 3464 0 -1 4610
box -4 -6 52 206
use OAI21X1  _4061_
timestamp 1596033377
transform 1 0 3464 0 -1 4610
box -4 -6 68 206
use AOI21X1  _4251_
timestamp 1596033377
transform -1 0 3592 0 -1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert292
timestamp 1596033377
transform 1 0 3592 0 -1 4610
box -4 -6 52 206
use AOI21X1  _4073_
timestamp 1596033377
transform -1 0 3704 0 -1 4610
box -4 -6 68 206
use OAI21X1  _2152_
timestamp 1596033377
transform -1 0 3768 0 -1 4610
box -4 -6 68 206
use INVX1  _2150_
timestamp 1596033377
transform -1 0 3800 0 -1 4610
box -4 -6 36 206
use NAND2X1  _2160_
timestamp 1596033377
transform 1 0 3800 0 -1 4610
box -4 -6 52 206
use OAI21X1  _2161_
timestamp 1596033377
transform -1 0 3912 0 -1 4610
box -4 -6 68 206
use OAI21X1  _2155_
timestamp 1596033377
transform 1 0 3912 0 -1 4610
box -4 -6 68 206
use NAND2X1  _2154_
timestamp 1596033377
transform 1 0 3976 0 -1 4610
box -4 -6 52 206
use DFFPOSX1  _4439_
timestamp 1596033377
transform -1 0 4216 0 -1 4610
box -4 -6 196 206
use DFFPOSX1  _4342_
timestamp 1596033377
transform 1 0 4216 0 -1 4610
box -4 -6 196 206
use FILL  SFILL44080x44100
timestamp 1596033377
transform -1 0 4424 0 -1 4610
box -4 -6 20 206
use NOR2X1  _3901_
timestamp 1596033377
transform -1 0 4520 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3902_
timestamp 1596033377
transform -1 0 4584 0 -1 4610
box -4 -6 68 206
use OAI21X1  _4010_
timestamp 1596033377
transform 1 0 4584 0 -1 4610
box -4 -6 68 206
use FILL  SFILL44240x44100
timestamp 1596033377
transform -1 0 4440 0 -1 4610
box -4 -6 20 206
use FILL  SFILL44400x44100
timestamp 1596033377
transform -1 0 4456 0 -1 4610
box -4 -6 20 206
use FILL  SFILL44560x44100
timestamp 1596033377
transform -1 0 4472 0 -1 4610
box -4 -6 20 206
use OAI22X1  _4011_
timestamp 1596033377
transform -1 0 4728 0 -1 4610
box -4 -6 84 206
use BUFX2  BUFX2_insert212
timestamp 1596033377
transform -1 0 4776 0 -1 4610
box -4 -6 52 206
use NOR2X1  _4009_
timestamp 1596033377
transform 1 0 4776 0 -1 4610
box -4 -6 52 206
use MUX2X1  _4249_
timestamp 1596033377
transform -1 0 4920 0 -1 4610
box -4 -6 100 206
use OAI22X1  _4248_
timestamp 1596033377
transform -1 0 5000 0 -1 4610
box -4 -6 84 206
use OAI21X1  _4247_
timestamp 1596033377
transform -1 0 5064 0 -1 4610
box -4 -6 68 206
use OAI21X1  _4069_
timestamp 1596033377
transform 1 0 5064 0 -1 4610
box -4 -6 68 206
use MUX2X1  _4067_
timestamp 1596033377
transform 1 0 5128 0 -1 4610
box -4 -6 100 206
use MUX2X1  _4245_
timestamp 1596033377
transform 1 0 5224 0 -1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert115
timestamp 1596033377
transform -1 0 5368 0 -1 4610
box -4 -6 52 206
use MUX2X1  _4179_
timestamp 1596033377
transform 1 0 5368 0 -1 4610
box -4 -6 100 206
use NOR2X1  _3676_
timestamp 1596033377
transform 1 0 5464 0 -1 4610
box -4 -6 52 206
use AOI21X1  _3677_
timestamp 1596033377
transform -1 0 5576 0 -1 4610
box -4 -6 68 206
use MUX2X1  _4001_
timestamp 1596033377
transform 1 0 5576 0 -1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert87
timestamp 1596033377
transform -1 0 5720 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert222
timestamp 1596033377
transform -1 0 5768 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert120
timestamp 1596033377
transform -1 0 5816 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert277
timestamp 1596033377
transform 1 0 5816 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert88
timestamp 1596033377
transform 1 0 5864 0 -1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert91
timestamp 1596033377
transform 1 0 5976 0 -1 4610
box -4 -6 52 206
use FILL  SFILL59120x44100
timestamp 1596033377
transform -1 0 5928 0 -1 4610
box -4 -6 20 206
use FILL  SFILL59280x44100
timestamp 1596033377
transform -1 0 5944 0 -1 4610
box -4 -6 20 206
use FILL  SFILL59440x44100
timestamp 1596033377
transform -1 0 5960 0 -1 4610
box -4 -6 20 206
use FILL  SFILL59600x44100
timestamp 1596033377
transform -1 0 5976 0 -1 4610
box -4 -6 20 206
use NOR2X1  _4235_
timestamp 1596033377
transform 1 0 6024 0 -1 4610
box -4 -6 52 206
use NOR2X1  _4053_
timestamp 1596033377
transform -1 0 6120 0 -1 4610
box -4 -6 52 206
use OAI22X1  _4055_
timestamp 1596033377
transform -1 0 6200 0 -1 4610
box -4 -6 84 206
use BUFX2  BUFX2_insert209
timestamp 1596033377
transform 1 0 6200 0 -1 4610
box -4 -6 52 206
use NOR2X1  _4231_
timestamp 1596033377
transform 1 0 6248 0 -1 4610
box -4 -6 52 206
use OAI21X1  _4054_
timestamp 1596033377
transform -1 0 6360 0 -1 4610
box -4 -6 68 206
use OAI22X1  _4233_
timestamp 1596033377
transform 1 0 6360 0 -1 4610
box -4 -6 84 206
use OAI21X1  _4232_
timestamp 1596033377
transform -1 0 6504 0 -1 4610
box -4 -6 68 206
use MUX2X1  _4230_
timestamp 1596033377
transform -1 0 6600 0 -1 4610
box -4 -6 100 206
use MUX2X1  _4052_
timestamp 1596033377
transform -1 0 6696 0 -1 4610
box -4 -6 100 206
use BUFX2  BUFX2_insert166
timestamp 1596033377
transform 1 0 6696 0 -1 4610
box -4 -6 52 206
use NOR2X1  _4280_
timestamp 1596033377
transform 1 0 6744 0 -1 4610
box -4 -6 52 206
use AOI21X1  _4281_
timestamp 1596033377
transform -1 0 6856 0 -1 4610
box -4 -6 68 206
use NOR2X1  _4290_
timestamp 1596033377
transform 1 0 6856 0 -1 4610
box -4 -6 52 206
use AOI21X1  _4291_
timestamp 1596033377
transform -1 0 6968 0 -1 4610
box -4 -6 68 206
use NOR2X1  _4292_
timestamp 1596033377
transform -1 0 7016 0 -1 4610
box -4 -6 52 206
use DFFPOSX1  _4422_
timestamp 1596033377
transform -1 0 7208 0 -1 4610
box -4 -6 196 206
use CLKBUF1  CLKBUF1_insert32
timestamp 1596033377
transform -1 0 7352 0 -1 4610
box -4 -6 148 206
use FILL  FILL70960x44100
timestamp 1596033377
transform -1 0 7368 0 -1 4610
box -4 -6 20 206
use FILL  FILL71120x44100
timestamp 1596033377
transform -1 0 7384 0 -1 4610
box -4 -6 20 206
use FILL  FILL71280x44100
timestamp 1596033377
transform -1 0 7400 0 -1 4610
box -4 -6 20 206
use AND2X2  _2520_
timestamp 1596033377
transform -1 0 72 0 1 4610
box -4 -6 68 206
use INVX1  _2518_
timestamp 1596033377
transform -1 0 104 0 1 4610
box -4 -6 36 206
use NOR2X1  _2519_
timestamp 1596033377
transform -1 0 152 0 1 4610
box -4 -6 52 206
use NAND2X1  _2516_
timestamp 1596033377
transform 1 0 152 0 1 4610
box -4 -6 52 206
use NOR2X1  _2242_
timestamp 1596033377
transform 1 0 200 0 1 4610
box -4 -6 52 206
use INVX1  _2240_
timestamp 1596033377
transform 1 0 248 0 1 4610
box -4 -6 36 206
use NOR2X1  _2243_
timestamp 1596033377
transform 1 0 280 0 1 4610
box -4 -6 52 206
use NOR2X1  _2241_
timestamp 1596033377
transform -1 0 376 0 1 4610
box -4 -6 52 206
use INVX1  _2239_
timestamp 1596033377
transform 1 0 376 0 1 4610
box -4 -6 36 206
use OAI21X1  _2253_
timestamp 1596033377
transform 1 0 408 0 1 4610
box -4 -6 68 206
use NAND2X1  _2249_
timestamp 1596033377
transform -1 0 520 0 1 4610
box -4 -6 52 206
use AND2X2  _2236_
timestamp 1596033377
transform -1 0 584 0 1 4610
box -4 -6 68 206
use NOR2X1  _2237_
timestamp 1596033377
transform 1 0 584 0 1 4610
box -4 -6 52 206
use AOI21X1  _2254_
timestamp 1596033377
transform -1 0 696 0 1 4610
box -4 -6 68 206
use INVX1  _2251_
timestamp 1596033377
transform -1 0 728 0 1 4610
box -4 -6 36 206
use INVX1  _2501_
timestamp 1596033377
transform 1 0 728 0 1 4610
box -4 -6 36 206
use NAND2X1  _2503_
timestamp 1596033377
transform -1 0 808 0 1 4610
box -4 -6 52 206
use INVX1  _2230_
timestamp 1596033377
transform 1 0 808 0 1 4610
box -4 -6 36 206
use OAI21X1  _2232_
timestamp 1596033377
transform -1 0 904 0 1 4610
box -4 -6 68 206
use NOR2X1  _2224_
timestamp 1596033377
transform -1 0 952 0 1 4610
box -4 -6 52 206
use NOR2X1  _2225_
timestamp 1596033377
transform 1 0 952 0 1 4610
box -4 -6 52 206
use OAI21X1  _2229_
timestamp 1596033377
transform 1 0 1000 0 1 4610
box -4 -6 68 206
use INVX1  _2222_
timestamp 1596033377
transform -1 0 1096 0 1 4610
box -4 -6 36 206
use OAI21X1  _2228_
timestamp 1596033377
transform 1 0 1096 0 1 4610
box -4 -6 68 206
use INVX1  _2217_
timestamp 1596033377
transform -1 0 1192 0 1 4610
box -4 -6 36 206
use NOR2X1  _2219_
timestamp 1596033377
transform -1 0 1240 0 1 4610
box -4 -6 52 206
use OAI21X1  _2221_
timestamp 1596033377
transform 1 0 1240 0 1 4610
box -4 -6 68 206
use NAND2X1  _2216_
timestamp 1596033377
transform -1 0 1352 0 1 4610
box -4 -6 52 206
use NOR2X1  _2218_
timestamp 1596033377
transform -1 0 1400 0 1 4610
box -4 -6 52 206
use FILL  SFILL14000x46100
timestamp 1596033377
transform 1 0 1400 0 1 4610
box -4 -6 20 206
use NAND2X1  _2592_
timestamp 1596033377
transform -1 0 1512 0 1 4610
box -4 -6 52 206
use AOI21X1  _2652_
timestamp 1596033377
transform 1 0 1512 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert173
timestamp 1596033377
transform -1 0 1624 0 1 4610
box -4 -6 52 206
use FILL  SFILL14160x46100
timestamp 1596033377
transform 1 0 1416 0 1 4610
box -4 -6 20 206
use FILL  SFILL14320x46100
timestamp 1596033377
transform 1 0 1432 0 1 4610
box -4 -6 20 206
use FILL  SFILL14480x46100
timestamp 1596033377
transform 1 0 1448 0 1 4610
box -4 -6 20 206
use XNOR2X1  _2574_
timestamp 1596033377
transform 1 0 1624 0 1 4610
box -4 -6 116 206
use NOR2X1  _2577_
timestamp 1596033377
transform -1 0 1784 0 1 4610
box -4 -6 52 206
use NAND2X1  _2576_
timestamp 1596033377
transform 1 0 1784 0 1 4610
box -4 -6 52 206
use XNOR2X1  _2575_
timestamp 1596033377
transform -1 0 1944 0 1 4610
box -4 -6 116 206
use BUFX2  BUFX2_insert107
timestamp 1596033377
transform 1 0 1944 0 1 4610
box -4 -6 52 206
use INVX1  _2854_
timestamp 1596033377
transform 1 0 1992 0 1 4610
box -4 -6 36 206
use AOI22X1  _2855_
timestamp 1596033377
transform -1 0 2104 0 1 4610
box -4 -6 84 206
use NAND3X1  _2860_
timestamp 1596033377
transform 1 0 2104 0 1 4610
box -4 -6 68 206
use OAI21X1  _2925_
timestamp 1596033377
transform -1 0 2232 0 1 4610
box -4 -6 68 206
use INVX1  _2853_
timestamp 1596033377
transform -1 0 2264 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert244
timestamp 1596033377
transform -1 0 2312 0 1 4610
box -4 -6 52 206
use AOI21X1  _2929_
timestamp 1596033377
transform 1 0 2312 0 1 4610
box -4 -6 68 206
use NOR2X1  _2861_
timestamp 1596033377
transform -1 0 2424 0 1 4610
box -4 -6 52 206
use NAND2X1  _2749_
timestamp 1596033377
transform -1 0 2472 0 1 4610
box -4 -6 52 206
use AND2X2  _2686_
timestamp 1596033377
transform 1 0 2472 0 1 4610
box -4 -6 68 206
use OAI21X1  _2928_
timestamp 1596033377
transform 1 0 2536 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert174
timestamp 1596033377
transform -1 0 2648 0 1 4610
box -4 -6 52 206
use NAND3X1  _2852_
timestamp 1596033377
transform -1 0 2712 0 1 4610
box -4 -6 68 206
use AOI21X1  _2926_
timestamp 1596033377
transform -1 0 2776 0 1 4610
box -4 -6 68 206
use INVX1  _2849_
timestamp 1596033377
transform 1 0 2776 0 1 4610
box -4 -6 36 206
use AOI22X1  _2851_
timestamp 1596033377
transform 1 0 2808 0 1 4610
box -4 -6 84 206
use INVX1  _2850_
timestamp 1596033377
transform -1 0 2920 0 1 4610
box -4 -6 36 206
use NAND2X1  _2846_
timestamp 1596033377
transform 1 0 2984 0 1 4610
box -4 -6 52 206
use FILL  SFILL29200x46100
timestamp 1596033377
transform 1 0 2920 0 1 4610
box -4 -6 20 206
use FILL  SFILL29360x46100
timestamp 1596033377
transform 1 0 2936 0 1 4610
box -4 -6 20 206
use FILL  SFILL29520x46100
timestamp 1596033377
transform 1 0 2952 0 1 4610
box -4 -6 20 206
use FILL  SFILL29680x46100
timestamp 1596033377
transform 1 0 2968 0 1 4610
box -4 -6 20 206
use INVX1  _2845_
timestamp 1596033377
transform -1 0 3064 0 1 4610
box -4 -6 36 206
use NAND2X1  _2668_
timestamp 1596033377
transform 1 0 3064 0 1 4610
box -4 -6 52 206
use INVX1  _2667_
timestamp 1596033377
transform -1 0 3144 0 1 4610
box -4 -6 36 206
use INVX1  _2141_
timestamp 1596033377
transform 1 0 3144 0 1 4610
box -4 -6 36 206
use BUFX2  BUFX2_insert193
timestamp 1596033377
transform -1 0 3224 0 1 4610
box -4 -6 52 206
use AND2X2  _2381_
timestamp 1596033377
transform -1 0 3288 0 1 4610
box -4 -6 68 206
use XNOR2X1  _2403_
timestamp 1596033377
transform 1 0 3288 0 1 4610
box -4 -6 116 206
use INVX1  _2147_
timestamp 1596033377
transform 1 0 3400 0 1 4610
box -4 -6 36 206
use INVX1  _2144_
timestamp 1596033377
transform 1 0 3432 0 1 4610
box -4 -6 36 206
use BUFX2  _2086_
timestamp 1596033377
transform -1 0 3512 0 1 4610
box -4 -6 52 206
use AOI21X1  _4062_
timestamp 1596033377
transform -1 0 3576 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4454_
timestamp 1596033377
transform -1 0 3768 0 1 4610
box -4 -6 196 206
use BUFX2  BUFX2_insert142
timestamp 1596033377
transform -1 0 3816 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert141
timestamp 1596033377
transform 1 0 3816 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4432_
timestamp 1596033377
transform -1 0 4056 0 1 4610
box -4 -6 196 206
use OAI21X1  _4184_
timestamp 1596033377
transform 1 0 4056 0 1 4610
box -4 -6 68 206
use AOI21X1  _4185_
timestamp 1596033377
transform -1 0 4184 0 1 4610
box -4 -6 68 206
use OAI21X1  _4261_
timestamp 1596033377
transform 1 0 4184 0 1 4610
box -4 -6 68 206
use OAI21X1  _4239_
timestamp 1596033377
transform -1 0 4312 0 1 4610
box -4 -6 68 206
use AOI21X1  _4262_
timestamp 1596033377
transform -1 0 4376 0 1 4610
box -4 -6 68 206
use FILL  SFILL43760x46100
timestamp 1596033377
transform 1 0 4376 0 1 4610
box -4 -6 20 206
use FILL  SFILL43920x46100
timestamp 1596033377
transform 1 0 4392 0 1 4610
box -4 -6 20 206
use FILL  SFILL44080x46100
timestamp 1596033377
transform 1 0 4408 0 1 4610
box -4 -6 20 206
use DFFPOSX1  _4321_
timestamp 1596033377
transform 1 0 4440 0 1 4610
box -4 -6 196 206
use FILL  SFILL44240x46100
timestamp 1596033377
transform 1 0 4424 0 1 4610
box -4 -6 20 206
use OAI21X1  _3758_
timestamp 1596033377
transform 1 0 4632 0 1 4610
box -4 -6 68 206
use NAND2X1  _3757_
timestamp 1596033377
transform -1 0 4744 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4369_
timestamp 1596033377
transform -1 0 4936 0 1 4610
box -4 -6 196 206
use OAI21X1  _3725_
timestamp 1596033377
transform 1 0 4936 0 1 4610
box -4 -6 68 206
use OAI21X1  _3724_
timestamp 1596033377
transform -1 0 5064 0 1 4610
box -4 -6 68 206
use NOR2X1  _4187_
timestamp 1596033377
transform 1 0 5064 0 1 4610
box -4 -6 52 206
use OAI22X1  _4189_
timestamp 1596033377
transform -1 0 5192 0 1 4610
box -4 -6 84 206
use OAI21X1  _4188_
timestamp 1596033377
transform 1 0 5192 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert12
timestamp 1596033377
transform -1 0 5304 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert282
timestamp 1596033377
transform -1 0 5352 0 1 4610
box -4 -6 52 206
use DFFPOSX1  _4400_
timestamp 1596033377
transform -1 0 5544 0 1 4610
box -4 -6 196 206
use OAI21X1  _3736_
timestamp 1596033377
transform -1 0 5608 0 1 4610
box -4 -6 68 206
use OAI21X1  _3726_
timestamp 1596033377
transform 1 0 5608 0 1 4610
box -4 -6 68 206
use OAI21X1  _3727_
timestamp 1596033377
transform -1 0 5736 0 1 4610
box -4 -6 68 206
use BUFX2  BUFX2_insert38
timestamp 1596033377
transform -1 0 5784 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert167
timestamp 1596033377
transform -1 0 5832 0 1 4610
box -4 -6 52 206
use BUFX2  BUFX2_insert281
timestamp 1596033377
transform 1 0 5832 0 1 4610
box -4 -6 52 206
use MUX2X1  _4060_
timestamp 1596033377
transform -1 0 5976 0 1 4610
box -4 -6 100 206
use FILL  SFILL59760x46100
timestamp 1596033377
transform 1 0 5976 0 1 4610
box -4 -6 20 206
use FILL  SFILL59920x46100
timestamp 1596033377
transform 1 0 5992 0 1 4610
box -4 -6 20 206
use FILL  SFILL60080x46100
timestamp 1596033377
transform 1 0 6008 0 1 4610
box -4 -6 20 206
use NOR2X1  _4057_
timestamp 1596033377
transform 1 0 6040 0 1 4610
box -4 -6 52 206
use OAI22X1  _4059_
timestamp 1596033377
transform 1 0 6088 0 1 4610
box -4 -6 84 206
use OAI21X1  _4058_
timestamp 1596033377
transform -1 0 6232 0 1 4610
box -4 -6 68 206
use FILL  SFILL60240x46100
timestamp 1596033377
transform 1 0 6024 0 1 4610
box -4 -6 20 206
use MUX2X1  _4238_
timestamp 1596033377
transform -1 0 6328 0 1 4610
box -4 -6 100 206
use OAI22X1  _4237_
timestamp 1596033377
transform 1 0 6328 0 1 4610
box -4 -6 84 206
use OAI21X1  _4236_
timestamp 1596033377
transform -1 0 6472 0 1 4610
box -4 -6 68 206
use NOR2X1  _3899_
timestamp 1596033377
transform 1 0 6472 0 1 4610
box -4 -6 52 206
use AOI21X1  _3900_
timestamp 1596033377
transform -1 0 6584 0 1 4610
box -4 -6 68 206
use DFFPOSX1  _4341_
timestamp 1596033377
transform -1 0 6776 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4416_
timestamp 1596033377
transform -1 0 6968 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4421_
timestamp 1596033377
transform -1 0 7160 0 1 4610
box -4 -6 196 206
use DFFPOSX1  _4389_
timestamp 1596033377
transform -1 0 7352 0 1 4610
box -4 -6 196 206
use FILL  FILL70960x46100
timestamp 1596033377
transform 1 0 7352 0 1 4610
box -4 -6 20 206
use FILL  FILL71120x46100
timestamp 1596033377
transform 1 0 7368 0 1 4610
box -4 -6 20 206
use FILL  FILL71280x46100
timestamp 1596033377
transform 1 0 7384 0 1 4610
box -4 -6 20 206
use XNOR2X1  _2582_
timestamp 1596033377
transform 1 0 8 0 -1 5010
box -4 -6 116 206
use OAI21X1  _2252_
timestamp 1596033377
transform 1 0 120 0 -1 5010
box -4 -6 68 206
use INVX1  _2515_
timestamp 1596033377
transform -1 0 216 0 -1 5010
box -4 -6 36 206
use NOR2X1  _2235_
timestamp 1596033377
transform -1 0 264 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert202
timestamp 1596033377
transform -1 0 312 0 -1 5010
box -4 -6 52 206
use BUFX2  _2102_
timestamp 1596033377
transform -1 0 360 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert161
timestamp 1596033377
transform -1 0 408 0 -1 5010
box -4 -6 52 206
use NOR2X1  _2591_
timestamp 1596033377
transform -1 0 456 0 -1 5010
box -4 -6 52 206
use NAND3X1  _2590_
timestamp 1596033377
transform -1 0 520 0 -1 5010
box -4 -6 68 206
use INVX1  _2588_
timestamp 1596033377
transform -1 0 552 0 -1 5010
box -4 -6 36 206
use AOI22X1  _2589_
timestamp 1596033377
transform 1 0 552 0 -1 5010
box -4 -6 84 206
use OR2X2  _2587_
timestamp 1596033377
transform -1 0 696 0 -1 5010
box -4 -6 68 206
use INVX1  _2586_
timestamp 1596033377
transform -1 0 728 0 -1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert229
timestamp 1596033377
transform -1 0 776 0 -1 5010
box -4 -6 52 206
use NOR2X1  _2320_
timestamp 1596033377
transform -1 0 824 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert80
timestamp 1596033377
transform -1 0 872 0 -1 5010
box -4 -6 52 206
use INVX1  _2223_
timestamp 1596033377
transform 1 0 872 0 -1 5010
box -4 -6 36 206
use INVX1  _2782_
timestamp 1596033377
transform 1 0 904 0 -1 5010
box -4 -6 36 206
use NAND2X1  _2783_
timestamp 1596033377
transform 1 0 936 0 -1 5010
box -4 -6 52 206
use OAI22X1  _2786_
timestamp 1596033377
transform -1 0 1064 0 -1 5010
box -4 -6 84 206
use BUFX2  BUFX2_insert44
timestamp 1596033377
transform -1 0 1112 0 -1 5010
box -4 -6 52 206
use INVX1  _2785_
timestamp 1596033377
transform -1 0 1144 0 -1 5010
box -4 -6 36 206
use AOI21X1  _2837_
timestamp 1596033377
transform 1 0 1144 0 -1 5010
box -4 -6 68 206
use INVX1  _2827_
timestamp 1596033377
transform -1 0 1240 0 -1 5010
box -4 -6 36 206
use OAI21X1  _2836_
timestamp 1596033377
transform -1 0 1304 0 -1 5010
box -4 -6 68 206
use NAND3X1  _2773_
timestamp 1596033377
transform 1 0 1304 0 -1 5010
box -4 -6 68 206
use OAI21X1  _2832_
timestamp 1596033377
transform -1 0 1432 0 -1 5010
box -4 -6 68 206
use INVX1  _2767_
timestamp 1596033377
transform -1 0 1528 0 -1 5010
box -4 -6 36 206
use INVX1  _2770_
timestamp 1596033377
transform 1 0 1528 0 -1 5010
box -4 -6 36 206
use AOI22X1  _2772_
timestamp 1596033377
transform 1 0 1560 0 -1 5010
box -4 -6 84 206
use FILL  SFILL14320x48100
timestamp 1596033377
transform -1 0 1448 0 -1 5010
box -4 -6 20 206
use FILL  SFILL14480x48100
timestamp 1596033377
transform -1 0 1464 0 -1 5010
box -4 -6 20 206
use FILL  SFILL14640x48100
timestamp 1596033377
transform -1 0 1480 0 -1 5010
box -4 -6 20 206
use FILL  SFILL14800x48100
timestamp 1596033377
transform -1 0 1496 0 -1 5010
box -4 -6 20 206
use INVX1  _2771_
timestamp 1596033377
transform -1 0 1672 0 -1 5010
box -4 -6 36 206
use INVX1  _2679_
timestamp 1596033377
transform 1 0 1672 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2681_
timestamp 1596033377
transform 1 0 1704 0 -1 5010
box -4 -6 84 206
use INVX1  _2680_
timestamp 1596033377
transform -1 0 1816 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2923_
timestamp 1596033377
transform 1 0 1816 0 -1 5010
box -4 -6 84 206
use OAI21X1  _2876_
timestamp 1596033377
transform 1 0 1896 0 -1 5010
box -4 -6 68 206
use NOR2X1  _2877_
timestamp 1596033377
transform -1 0 2008 0 -1 5010
box -4 -6 52 206
use NAND3X1  _2869_
timestamp 1596033377
transform -1 0 2072 0 -1 5010
box -4 -6 68 206
use INVX1  _2683_
timestamp 1596033377
transform 1 0 2072 0 -1 5010
box -4 -6 36 206
use OAI22X1  _2684_
timestamp 1596033377
transform -1 0 2184 0 -1 5010
box -4 -6 84 206
use NOR2X1  _2685_
timestamp 1596033377
transform -1 0 2232 0 -1 5010
box -4 -6 52 206
use INVX1  _2682_
timestamp 1596033377
transform -1 0 2264 0 -1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert76
timestamp 1596033377
transform 1 0 2264 0 -1 5010
box -4 -6 52 206
use AOI21X1  _2835_
timestamp 1596033377
transform -1 0 2376 0 -1 5010
box -4 -6 68 206
use INVX1  _2763_
timestamp 1596033377
transform 1 0 2376 0 -1 5010
box -4 -6 36 206
use NOR2X1  _2766_
timestamp 1596033377
transform 1 0 2408 0 -1 5010
box -4 -6 52 206
use OAI22X1  _2765_
timestamp 1596033377
transform 1 0 2456 0 -1 5010
box -4 -6 84 206
use NAND2X1  _2833_
timestamp 1596033377
transform -1 0 2584 0 -1 5010
box -4 -6 52 206
use INVX1  _2764_
timestamp 1596033377
transform -1 0 2616 0 -1 5010
box -4 -6 36 206
use NAND2X1  _2868_
timestamp 1596033377
transform 1 0 2616 0 -1 5010
box -4 -6 52 206
use INVX1  _2867_
timestamp 1596033377
transform -1 0 2696 0 -1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert99
timestamp 1596033377
transform 1 0 2696 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert233
timestamp 1596033377
transform -1 0 2792 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert204
timestamp 1596033377
transform 1 0 2792 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert159
timestamp 1596033377
transform 1 0 2840 0 -1 5010
box -4 -6 52 206
use NAND2X1  _2145_
timestamp 1596033377
transform 1 0 2888 0 -1 5010
box -4 -6 52 206
use OAI21X1  _2146_
timestamp 1596033377
transform -1 0 3064 0 -1 5010
box -4 -6 68 206
use FILL  SFILL29360x48100
timestamp 1596033377
transform -1 0 2952 0 -1 5010
box -4 -6 20 206
use FILL  SFILL29520x48100
timestamp 1596033377
transform -1 0 2968 0 -1 5010
box -4 -6 20 206
use FILL  SFILL29680x48100
timestamp 1596033377
transform -1 0 2984 0 -1 5010
box -4 -6 20 206
use FILL  SFILL29840x48100
timestamp 1596033377
transform -1 0 3000 0 -1 5010
box -4 -6 20 206
use OAI21X1  _2143_
timestamp 1596033377
transform 1 0 3064 0 -1 5010
box -4 -6 68 206
use NAND2X1  _2142_
timestamp 1596033377
transform 1 0 3128 0 -1 5010
box -4 -6 52 206
use OAI21X1  _4006_
timestamp 1596033377
transform 1 0 3176 0 -1 5010
box -4 -6 68 206
use AOI21X1  _4007_
timestamp 1596033377
transform -1 0 3304 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4039_
timestamp 1596033377
transform 1 0 3304 0 -1 5010
box -4 -6 68 206
use AOI21X1  _4040_
timestamp 1596033377
transform -1 0 3432 0 -1 5010
box -4 -6 68 206
use BUFX2  _2090_
timestamp 1596033377
transform -1 0 3480 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert77
timestamp 1596033377
transform -1 0 3528 0 -1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert140
timestamp 1596033377
transform -1 0 3576 0 -1 5010
box -4 -6 52 206
use OAI21X1  _4083_
timestamp 1596033377
transform 1 0 3576 0 -1 5010
box -4 -6 68 206
use AOI21X1  _4084_
timestamp 1596033377
transform -1 0 3704 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4455_
timestamp 1596033377
transform -1 0 3896 0 -1 5010
box -4 -6 196 206
use OAI21X1  _4195_
timestamp 1596033377
transform -1 0 3960 0 -1 5010
box -4 -6 68 206
use AOI21X1  _4196_
timestamp 1596033377
transform -1 0 4024 0 -1 5010
box -4 -6 68 206
use INVX4  _3696_
timestamp 1596033377
transform -1 0 4072 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4306_
timestamp 1596033377
transform 1 0 4072 0 -1 5010
box -4 -6 196 206
use AOI21X1  _4240_
timestamp 1596033377
transform -1 0 4328 0 -1 5010
box -4 -6 68 206
use AOI21X1  _3892_
timestamp 1596033377
transform 1 0 4328 0 -1 5010
box -4 -6 68 206
use NOR2X1  _3891_
timestamp 1596033377
transform -1 0 4440 0 -1 5010
box -4 -6 52 206
use NAND2X1  _3860_
timestamp 1596033377
transform 1 0 4504 0 -1 5010
box -4 -6 52 206
use OAI21X1  _3861_
timestamp 1596033377
transform -1 0 4616 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4014_
timestamp 1596033377
transform 1 0 4616 0 -1 5010
box -4 -6 68 206
use FILL  SFILL44400x48100
timestamp 1596033377
transform -1 0 4456 0 -1 5010
box -4 -6 20 206
use FILL  SFILL44560x48100
timestamp 1596033377
transform -1 0 4472 0 -1 5010
box -4 -6 20 206
use FILL  SFILL44720x48100
timestamp 1596033377
transform -1 0 4488 0 -1 5010
box -4 -6 20 206
use FILL  SFILL44880x48100
timestamp 1596033377
transform -1 0 4504 0 -1 5010
box -4 -6 20 206
use OAI21X1  _4192_
timestamp 1596033377
transform 1 0 4680 0 -1 5010
box -4 -6 68 206
use MUX2X1  _4194_
timestamp 1596033377
transform -1 0 4840 0 -1 5010
box -4 -6 100 206
use DFFPOSX1  _4338_
timestamp 1596033377
transform 1 0 4840 0 -1 5010
box -4 -6 196 206
use NOR2X1  _3893_
timestamp 1596033377
transform -1 0 5080 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3894_
timestamp 1596033377
transform -1 0 5144 0 -1 5010
box -4 -6 68 206
use MUX2X1  _4260_
timestamp 1596033377
transform -1 0 5240 0 -1 5010
box -4 -6 100 206
use DFFPOSX1  _4375_
timestamp 1596033377
transform 1 0 5240 0 -1 5010
box -4 -6 196 206
use OAI21X1  _3737_
timestamp 1596033377
transform 1 0 5432 0 -1 5010
box -4 -6 68 206
use DFFPOSX1  _4370_
timestamp 1596033377
transform 1 0 5496 0 -1 5010
box -4 -6 196 206
use NOR2X1  _4075_
timestamp 1596033377
transform 1 0 5688 0 -1 5010
box -4 -6 52 206
use OAI22X1  _4077_
timestamp 1596033377
transform 1 0 5736 0 -1 5010
box -4 -6 84 206
use MUX2X1  _4082_
timestamp 1596033377
transform 1 0 5816 0 -1 5010
box -4 -6 100 206
use NOR2X1  _4257_
timestamp 1596033377
transform -1 0 6024 0 -1 5010
box -4 -6 52 206
use FILL  SFILL59120x48100
timestamp 1596033377
transform -1 0 5928 0 -1 5010
box -4 -6 20 206
use FILL  SFILL59280x48100
timestamp 1596033377
transform -1 0 5944 0 -1 5010
box -4 -6 20 206
use FILL  SFILL59440x48100
timestamp 1596033377
transform -1 0 5960 0 -1 5010
box -4 -6 20 206
use FILL  SFILL59600x48100
timestamp 1596033377
transform -1 0 5976 0 -1 5010
box -4 -6 20 206
use OAI22X1  _4259_
timestamp 1596033377
transform 1 0 6024 0 -1 5010
box -4 -6 84 206
use NOR2X1  _4079_
timestamp 1596033377
transform -1 0 6152 0 -1 5010
box -4 -6 52 206
use OAI22X1  _4081_
timestamp 1596033377
transform 1 0 6152 0 -1 5010
box -4 -6 84 206
use OAI21X1  _4080_
timestamp 1596033377
transform -1 0 6296 0 -1 5010
box -4 -6 68 206
use OAI21X1  _4258_
timestamp 1596033377
transform -1 0 6360 0 -1 5010
box -4 -6 68 206
use MUX2X1  _4256_
timestamp 1596033377
transform -1 0 6456 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4078_
timestamp 1596033377
transform -1 0 6552 0 -1 5010
box -4 -6 100 206
use NOR2X1  _3903_
timestamp 1596033377
transform 1 0 6552 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3904_
timestamp 1596033377
transform 1 0 6600 0 -1 5010
box -4 -6 68 206
use MUX2X1  _4234_
timestamp 1596033377
transform 1 0 6664 0 -1 5010
box -4 -6 100 206
use MUX2X1  _4056_
timestamp 1596033377
transform 1 0 6760 0 -1 5010
box -4 -6 100 206
use BUFX2  BUFX2_insert220
timestamp 1596033377
transform 1 0 6856 0 -1 5010
box -4 -6 52 206
use NOR2X1  _3697_
timestamp 1596033377
transform -1 0 6952 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3698_
timestamp 1596033377
transform -1 0 7016 0 -1 5010
box -4 -6 68 206
use NOR2X1  _3691_
timestamp 1596033377
transform -1 0 7064 0 -1 5010
box -4 -6 52 206
use AOI21X1  _3692_
timestamp 1596033377
transform -1 0 7128 0 -1 5010
box -4 -6 68 206
use NAND2X1  _3799_
timestamp 1596033377
transform -1 0 7176 0 -1 5010
box -4 -6 52 206
use DFFPOSX1  _4407_
timestamp 1596033377
transform -1 0 7368 0 -1 5010
box -4 -6 196 206
use FILL  FILL71120x48100
timestamp 1596033377
transform -1 0 7384 0 -1 5010
box -4 -6 20 206
use FILL  FILL71280x48100
timestamp 1596033377
transform -1 0 7400 0 -1 5010
box -4 -6 20 206
use XNOR2X1  _2511_
timestamp 1596033377
transform 1 0 8 0 1 5010
box -4 -6 116 206
use AND2X2  _2233_
timestamp 1596033377
transform 1 0 120 0 1 5010
box -4 -6 68 206
use NOR2X1  _2234_
timestamp 1596033377
transform -1 0 232 0 1 5010
box -4 -6 52 206
use INVX1  _2580_
timestamp 1596033377
transform 1 0 232 0 1 5010
box -4 -6 36 206
use NAND2X1  _2581_
timestamp 1596033377
transform -1 0 312 0 1 5010
box -4 -6 52 206
use NAND3X1  _2583_
timestamp 1596033377
transform 1 0 312 0 1 5010
box -4 -6 68 206
use NAND3X1  _2641_
timestamp 1596033377
transform 1 0 376 0 1 5010
box -4 -6 68 206
use OAI22X1  _2642_
timestamp 1596033377
transform 1 0 440 0 1 5010
box -4 -6 84 206
use AOI22X1  _2640_
timestamp 1596033377
transform 1 0 520 0 1 5010
box -4 -6 84 206
use NAND2X1  _2585_
timestamp 1596033377
transform -1 0 648 0 1 5010
box -4 -6 52 206
use INVX1  _2584_
timestamp 1596033377
transform -1 0 680 0 1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert160
timestamp 1596033377
transform 1 0 680 0 1 5010
box -4 -6 52 206
use AND2X2  _2319_
timestamp 1596033377
transform 1 0 728 0 1 5010
box -4 -6 68 206
use NOR2X1  _2318_
timestamp 1596033377
transform -1 0 840 0 1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert79
timestamp 1596033377
transform -1 0 888 0 1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert230
timestamp 1596033377
transform -1 0 936 0 1 5010
box -4 -6 52 206
use OAI21X1  _2831_
timestamp 1596033377
transform 1 0 936 0 1 5010
box -4 -6 68 206
use OAI21X1  _2830_
timestamp 1596033377
transform 1 0 1000 0 1 5010
box -4 -6 68 206
use NOR2X1  _2787_
timestamp 1596033377
transform 1 0 1064 0 1 5010
box -4 -6 52 206
use NAND2X1  _2788_
timestamp 1596033377
transform 1 0 1112 0 1 5010
box -4 -6 52 206
use OAI21X1  _2784_
timestamp 1596033377
transform -1 0 1224 0 1 5010
box -4 -6 68 206
use NOR2X1  _2789_
timestamp 1596033377
transform -1 0 1272 0 1 5010
box -4 -6 52 206
use INVX1  _2781_
timestamp 1596033377
transform -1 0 1304 0 1 5010
box -4 -6 36 206
use BUFX2  BUFX2_insert231
timestamp 1596033377
transform 1 0 1304 0 1 5010
box -4 -6 52 206
use AND2X2  _2366_
timestamp 1596033377
transform 1 0 1352 0 1 5010
box -4 -6 68 206
use AOI22X1  _2769_
timestamp 1596033377
transform 1 0 1480 0 1 5010
box -4 -6 84 206
use INVX1  _2768_
timestamp 1596033377
transform -1 0 1592 0 1 5010
box -4 -6 36 206
use NOR2X1  _2921_
timestamp 1596033377
transform -1 0 1640 0 1 5010
box -4 -6 52 206
use FILL  SFILL14160x50100
timestamp 1596033377
transform 1 0 1416 0 1 5010
box -4 -6 20 206
use FILL  SFILL14320x50100
timestamp 1596033377
transform 1 0 1432 0 1 5010
box -4 -6 20 206
use FILL  SFILL14480x50100
timestamp 1596033377
transform 1 0 1448 0 1 5010
box -4 -6 20 206
use FILL  SFILL14640x50100
timestamp 1596033377
transform 1 0 1464 0 1 5010
box -4 -6 20 206
use BUFX2  BUFX2_insert78
timestamp 1596033377
transform 1 0 1640 0 1 5010
box -4 -6 52 206
use INVX1  _2871_
timestamp 1596033377
transform 1 0 1688 0 1 5010
box -4 -6 36 206
use OAI22X1  _2873_
timestamp 1596033377
transform 1 0 1720 0 1 5010
box -4 -6 84 206
use INVX1  _2874_
timestamp 1596033377
transform 1 0 1800 0 1 5010
box -4 -6 36 206
use INVX1  _2872_
timestamp 1596033377
transform -1 0 1864 0 1 5010
box -4 -6 36 206
use OAI21X1  _2922_
timestamp 1596033377
transform -1 0 1928 0 1 5010
box -4 -6 68 206
use NAND2X1  _2875_
timestamp 1596033377
transform -1 0 1976 0 1 5010
box -4 -6 52 206
use INVX1  _2865_
timestamp 1596033377
transform 1 0 1976 0 1 5010
box -4 -6 36 206
use NAND2X1  _2866_
timestamp 1596033377
transform -1 0 2056 0 1 5010
box -4 -6 52 206
use NOR2X1  _2678_
timestamp 1596033377
transform -1 0 2104 0 1 5010
box -4 -6 52 206
use OAI21X1  _2736_
timestamp 1596033377
transform 1 0 2104 0 1 5010
box -4 -6 68 206
use OAI21X1  _2735_
timestamp 1596033377
transform -1 0 2232 0 1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert162
timestamp 1596033377
transform 1 0 2232 0 1 5010
box -4 -6 52 206
use AOI21X1  _2834_
timestamp 1596033377
transform 1 0 2280 0 1 5010
box -4 -6 68 206
use INVX1  _2760_
timestamp 1596033377
transform -1 0 2376 0 1 5010
box -4 -6 36 206
use OAI22X1  _2762_
timestamp 1596033377
transform 1 0 2376 0 1 5010
box -4 -6 84 206
use INVX1  _2761_
timestamp 1596033377
transform -1 0 2488 0 1 5010
box -4 -6 36 206
use BUFX2  _2111_
timestamp 1596033377
transform 1 0 2488 0 1 5010
box -4 -6 52 206
use BUFX2  BUFX2_insert43
timestamp 1596033377
transform -1 0 2584 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4448_
timestamp 1596033377
transform -1 0 2776 0 1 5010
box -4 -6 196 206
use NAND2X1  _2148_
timestamp 1596033377
transform -1 0 2824 0 1 5010
box -4 -6 52 206
use OAI21X1  _2149_
timestamp 1596033377
transform -1 0 2888 0 1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert232
timestamp 1596033377
transform 1 0 2888 0 1 5010
box -4 -6 52 206
use BUFX2  _2095_
timestamp 1596033377
transform -1 0 3048 0 1 5010
box -4 -6 52 206
use FILL  SFILL29360x50100
timestamp 1596033377
transform 1 0 2936 0 1 5010
box -4 -6 20 206
use FILL  SFILL29520x50100
timestamp 1596033377
transform 1 0 2952 0 1 5010
box -4 -6 20 206
use FILL  SFILL29680x50100
timestamp 1596033377
transform 1 0 2968 0 1 5010
box -4 -6 20 206
use FILL  SFILL29840x50100
timestamp 1596033377
transform 1 0 2984 0 1 5010
box -4 -6 20 206
use DFFPOSX1  _4435_
timestamp 1596033377
transform -1 0 3240 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4449_
timestamp 1596033377
transform -1 0 3432 0 1 5010
box -4 -6 196 206
use OAI21X1  _4017_
timestamp 1596033377
transform 1 0 3432 0 1 5010
box -4 -6 68 206
use AOI21X1  _4018_
timestamp 1596033377
transform -1 0 3560 0 1 5010
box -4 -6 68 206
use BUFX2  BUFX2_insert291
timestamp 1596033377
transform 1 0 3560 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4433_
timestamp 1596033377
transform -1 0 3800 0 1 5010
box -4 -6 196 206
use BUFX2  _2087_
timestamp 1596033377
transform -1 0 3848 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4437_
timestamp 1596033377
transform -1 0 4040 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4305_
timestamp 1596033377
transform 1 0 4040 0 1 5010
box -4 -6 196 206
use OAI21X1  _3859_
timestamp 1596033377
transform 1 0 4232 0 1 5010
box -4 -6 68 206
use NAND2X1  _3858_
timestamp 1596033377
transform -1 0 4344 0 1 5010
box -4 -6 52 206
use DFFPOSX1  _4337_
timestamp 1596033377
transform 1 0 4408 0 1 5010
box -4 -6 196 206
use FILL  SFILL43440x50100
timestamp 1596033377
transform 1 0 4344 0 1 5010
box -4 -6 20 206
use FILL  SFILL43600x50100
timestamp 1596033377
transform 1 0 4360 0 1 5010
box -4 -6 20 206
use FILL  SFILL43760x50100
timestamp 1596033377
transform 1 0 4376 0 1 5010
box -4 -6 20 206
use FILL  SFILL43920x50100
timestamp 1596033377
transform 1 0 4392 0 1 5010
box -4 -6 20 206
use OAI22X1  _4015_
timestamp 1596033377
transform -1 0 4680 0 1 5010
box -4 -6 84 206
use MUX2X1  _4016_
timestamp 1596033377
transform -1 0 4776 0 1 5010
box -4 -6 100 206
use OAI22X1  _4193_
timestamp 1596033377
transform -1 0 4856 0 1 5010
box -4 -6 84 206
use NOR2X1  _4013_
timestamp 1596033377
transform 1 0 4856 0 1 5010
box -4 -6 52 206
use NOR2X1  _4191_
timestamp 1596033377
transform 1 0 4904 0 1 5010
box -4 -6 52 206
use NOR2X1  _4202_
timestamp 1596033377
transform -1 0 5000 0 1 5010
box -4 -6 52 206
use OAI22X1  _4204_
timestamp 1596033377
transform 1 0 5000 0 1 5010
box -4 -6 84 206
use OAI21X1  _4203_
timestamp 1596033377
transform -1 0 5144 0 1 5010
box -4 -6 68 206
use NOR2X1  _4024_
timestamp 1596033377
transform -1 0 5192 0 1 5010
box -4 -6 52 206
use OAI21X1  _4025_
timestamp 1596033377
transform 1 0 5192 0 1 5010
box -4 -6 68 206
use OAI22X1  _4026_
timestamp 1596033377
transform 1 0 5256 0 1 5010
box -4 -6 84 206
use MUX2X1  _4027_
timestamp 1596033377
transform -1 0 5432 0 1 5010
box -4 -6 100 206
use OAI21X1  _4076_
timestamp 1596033377
transform -1 0 5496 0 1 5010
box -4 -6 68 206
use OAI21X1  _4254_
timestamp 1596033377
transform 1 0 5496 0 1 5010
box -4 -6 68 206
use OAI22X1  _4255_
timestamp 1596033377
transform -1 0 5640 0 1 5010
box -4 -6 84 206
use NOR2X1  _4253_
timestamp 1596033377
transform 1 0 5640 0 1 5010
box -4 -6 52 206
use NOR2X1  _4198_
timestamp 1596033377
transform -1 0 5736 0 1 5010
box -4 -6 52 206
use NOR2X1  _4020_
timestamp 1596033377
transform 1 0 5736 0 1 5010
box -4 -6 52 206
use OAI22X1  _4022_
timestamp 1596033377
transform 1 0 5784 0 1 5010
box -4 -6 84 206
use OAI21X1  _4021_
timestamp 1596033377
transform 1 0 5864 0 1 5010
box -4 -6 68 206
use MUX2X1  _4201_
timestamp 1596033377
transform 1 0 5992 0 1 5010
box -4 -6 100 206
use FILL  SFILL59280x50100
timestamp 1596033377
transform 1 0 5928 0 1 5010
box -4 -6 20 206
use FILL  SFILL59440x50100
timestamp 1596033377
transform 1 0 5944 0 1 5010
box -4 -6 20 206
use FILL  SFILL59600x50100
timestamp 1596033377
transform 1 0 5960 0 1 5010
box -4 -6 20 206
use FILL  SFILL59760x50100
timestamp 1596033377
transform 1 0 5976 0 1 5010
box -4 -6 20 206
use MUX2X1  _4023_
timestamp 1596033377
transform -1 0 6184 0 1 5010
box -4 -6 100 206
use NOR2X1  _4284_
timestamp 1596033377
transform -1 0 6232 0 1 5010
box -4 -6 52 206
use AOI21X1  _4285_
timestamp 1596033377
transform -1 0 6296 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4418_
timestamp 1596033377
transform -1 0 6488 0 1 5010
box -4 -6 196 206
use NOR2X1  _4294_
timestamp 1596033377
transform 1 0 6488 0 1 5010
box -4 -6 52 206
use AOI21X1  _4295_
timestamp 1596033377
transform -1 0 6600 0 1 5010
box -4 -6 68 206
use DFFPOSX1  _4423_
timestamp 1596033377
transform -1 0 6792 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4343_
timestamp 1596033377
transform -1 0 6984 0 1 5010
box -4 -6 196 206
use DFFPOSX1  _4402_
timestamp 1596033377
transform -1 0 7176 0 1 5010
box -4 -6 196 206
use NOR2X1  _3682_
timestamp 1596033377
transform 1 0 7176 0 1 5010
box -4 -6 52 206
use AOI21X1  _3683_
timestamp 1596033377
transform -1 0 7288 0 1 5010
box -4 -6 68 206
use OAI21X1  _3740_
timestamp 1596033377
transform 1 0 7288 0 1 5010
box -4 -6 68 206
use FILL  FILL70960x50100
timestamp 1596033377
transform 1 0 7352 0 1 5010
box -4 -6 20 206
use FILL  FILL71120x50100
timestamp 1596033377
transform 1 0 7368 0 1 5010
box -4 -6 20 206
use FILL  FILL71280x50100
timestamp 1596033377
transform 1 0 7384 0 1 5010
box -4 -6 20 206
use BUFX2  _2098_
timestamp 1596033377
transform -1 0 56 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert252
timestamp 1596033377
transform -1 0 104 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert254
timestamp 1596033377
transform 1 0 104 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert15
timestamp 1596033377
transform -1 0 200 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert17
timestamp 1596033377
transform 1 0 200 0 -1 5410
box -4 -6 52 206
use INVX1  _2578_
timestamp 1596033377
transform 1 0 248 0 -1 5410
box -4 -6 36 206
use NAND2X1  _2579_
timestamp 1596033377
transform -1 0 328 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert205
timestamp 1596033377
transform 1 0 328 0 -1 5410
box -4 -6 52 206
use AOI22X1  _2637_
timestamp 1596033377
transform -1 0 456 0 -1 5410
box -4 -6 84 206
use NOR2X1  _2638_
timestamp 1596033377
transform -1 0 504 0 -1 5410
box -4 -6 52 206
use INVX1  _2636_
timestamp 1596033377
transform -1 0 536 0 -1 5410
box -4 -6 36 206
use INVX1  _2639_
timestamp 1596033377
transform 1 0 536 0 -1 5410
box -4 -6 36 206
use BUFX2  _2099_
timestamp 1596033377
transform 1 0 568 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert16
timestamp 1596033377
transform -1 0 664 0 -1 5410
box -4 -6 52 206
use NAND2X1  _2778_
timestamp 1596033377
transform 1 0 664 0 -1 5410
box -4 -6 52 206
use OAI21X1  _2779_
timestamp 1596033377
transform -1 0 776 0 -1 5410
box -4 -6 68 206
use INVX1  _2775_
timestamp 1596033377
transform -1 0 808 0 -1 5410
box -4 -6 36 206
use INVX1  _2777_
timestamp 1596033377
transform 1 0 808 0 -1 5410
box -4 -6 36 206
use NOR2X1  _2780_
timestamp 1596033377
transform -1 0 888 0 -1 5410
box -4 -6 52 206
use OR2X2  _2828_
timestamp 1596033377
transform 1 0 888 0 -1 5410
box -4 -6 68 206
use OAI21X1  _2829_
timestamp 1596033377
transform 1 0 952 0 -1 5410
box -4 -6 68 206
use OAI22X1  _2776_
timestamp 1596033377
transform 1 0 1016 0 -1 5410
box -4 -6 84 206
use INVX1  _2774_
timestamp 1596033377
transform -1 0 1128 0 -1 5410
box -4 -6 36 206
use BUFX2  BUFX2_insert201
timestamp 1596033377
transform -1 0 1176 0 -1 5410
box -4 -6 52 206
use BUFX2  BUFX2_insert253
timestamp 1596033377
transform 1 0 1176 0 -1 5410
box -4 -6 52 206
use BUFX2  _2101_
timestamp 1596033377
transform 1 0 1224 0 -1 5410
box -4 -6 52 206
use INVX1  _2863_
timestamp 1596033377
transform 1 0 1272 0 -1 5410
box -4 -6 36 206
use AOI22X1  _2864_
timestamp 1596033377
transform -1 0 1384 0 -1 5410
box -4 -6 84 206
use INVX1  _2862_
timestamp 1596033377
transform -1 0 1416 0 -1 5410
box -4 -6 36 206
use INVX1  _2673_
timestamp 1596033377
transform 1 0 1480 0 -1 5410
box -4 -6 36 206
use BUFX2  _2100_
timestamp 1596033377
transform 1 0 1512 0 -1 5410
box -4 -6 52 206
use NAND2X1  _2732_
timestamp 1596033377
transform 1 0 1560 0 -1 5410
box -4 -6 52 206
use INVX1  _2672_
timestamp 1596033377
transform 1 0 1608 0 -1 5410
box -4 -6 36 206
use FILL  SFILL14160x52100
timestamp 1596033377
transform -1 0 1432 0 -1 5410
box -4 -6 20 206
use FILL  SFILL14320x52100
timestamp 1596033377
transform -1 0 1448 0 -1 5410
box -4 -6 20 206
use FILL  SFILL14480x52100
timestamp 1596033377
transform -1 0 1464 0 -1 5410
box -4 -6 20 206
use FILL  SFILL14640x52100
timestamp 1596033377
transform -1 0 1480 0 -1 5410
box -4 -6 20 206
use OAI22X1  _2674_
timestamp 1596033377
transform -1 0 1720 0 -1 5410
box -4 -6 84 206
use NAND2X1  _2731_
timestamp 1596033377
transform -1 0 1768 0 -1 5410
box -4 -6 52 206
use NAND3X1  _2733_
timestamp 1596033377
transform 1 0 1768 0 -1 5410
box -4 -6 68 206
use INVX1  _2676_
timestamp 1596033377
transform 1 0 1832 0 -1 5410
box -4 -6 36 206
use BUFX2  BUFX2_insert203
timestamp 1596033377
transform 1 0 1864 0 -1 5410
box -4 -6 52 206
use AOI22X1  _2730_
timestamp 1596033377
transform -1 0 1992 0 -1 5410
box -4 -6 84 206
use INVX1  _2675_
timestamp 1596033377
transform -1 0 2024 0 -1 5410
box -4 -6 36 206
use OAI22X1  _2677_
timestamp 1596033377
transform -1 0 2104 0 -1 5410
box -4 -6 84 206
use OAI21X1  _2734_
timestamp 1596033377
transform 1 0 2104 0 -1 5410
box -4 -6 68 206
use BUFX2  BUFX2_insert14
timestamp 1596033377
transform 1 0 2168 0 -1 5410
box -4 -6 52 206
use XOR2X1  _2374_
timestamp 1596033377
transform 1 0 2216 0 -1 5410
box -4 -6 116 206
use NOR2X1  _2376_
timestamp 1596033377
transform 1 0 2328 0 -1 5410
box -4 -6 52 206
use XOR2X1  _2375_
timestamp 1596033377
transform 1 0 2376 0 -1 5410
box -4 -6 116 206
use BUFX2  BUFX2_insert251
timestamp 1596033377
transform -1 0 2536 0 -1 5410
box -4 -6 52 206
use BUFX2  _2110_
timestamp 1596033377
transform 1 0 2536 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4434_
timestamp 1596033377
transform -1 0 2776 0 -1 5410
box -4 -6 196 206
use BUFX2  _2082_
timestamp 1596033377
transform 1 0 2776 0 -1 5410
box -4 -6 52 206
use BUFX2  _2083_
timestamp 1596033377
transform 1 0 2824 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4450_
timestamp 1596033377
transform -1 0 3128 0 -1 5410
box -4 -6 196 206
use FILL  SFILL28720x52100
timestamp 1596033377
transform -1 0 2888 0 -1 5410
box -4 -6 20 206
use FILL  SFILL28880x52100
timestamp 1596033377
transform -1 0 2904 0 -1 5410
box -4 -6 20 206
use FILL  SFILL29040x52100
timestamp 1596033377
transform -1 0 2920 0 -1 5410
box -4 -6 20 206
use FILL  SFILL29200x52100
timestamp 1596033377
transform -1 0 2936 0 -1 5410
box -4 -6 20 206
use DFFPOSX1  _4451_
timestamp 1596033377
transform -1 0 3320 0 -1 5410
box -4 -6 196 206
use OAI21X1  _4028_
timestamp 1596033377
transform 1 0 3320 0 -1 5410
box -4 -6 68 206
use AOI21X1  _4029_
timestamp 1596033377
transform -1 0 3448 0 -1 5410
box -4 -6 68 206
use OAI21X1  _4206_
timestamp 1596033377
transform 1 0 3448 0 -1 5410
box -4 -6 68 206
use AOI21X1  _4207_
timestamp 1596033377
transform -1 0 3576 0 -1 5410
box -4 -6 68 206
use BUFX2  _2103_
timestamp 1596033377
transform 1 0 3576 0 -1 5410
box -4 -6 52 206
use BUFX2  _2084_
timestamp 1596033377
transform 1 0 3624 0 -1 5410
box -4 -6 52 206
use BUFX2  _2085_
timestamp 1596033377
transform 1 0 3672 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4401_
timestamp 1596033377
transform -1 0 3912 0 -1 5410
box -4 -6 196 206
use NOR2X1  _3679_
timestamp 1596033377
transform 1 0 3912 0 -1 5410
box -4 -6 52 206
use AOI21X1  _3680_
timestamp 1596033377
transform -1 0 4024 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4311_
timestamp 1596033377
transform 1 0 4024 0 -1 5410
box -4 -6 196 206
use OAI21X1  _3871_
timestamp 1596033377
transform 1 0 4216 0 -1 5410
box -4 -6 68 206
use NAND2X1  _3870_
timestamp 1596033377
transform -1 0 4328 0 -1 5410
box -4 -6 52 206
use MUX2X1  _4012_
timestamp 1596033377
transform -1 0 4424 0 -1 5410
box -4 -6 100 206
use MUX2X1  _4190_
timestamp 1596033377
transform -1 0 4584 0 -1 5410
box -4 -6 100 206
use NOR2X1  _4282_
timestamp 1596033377
transform 1 0 4584 0 -1 5410
box -4 -6 52 206
use FILL  SFILL44240x52100
timestamp 1596033377
transform -1 0 4440 0 -1 5410
box -4 -6 20 206
use FILL  SFILL44400x52100
timestamp 1596033377
transform -1 0 4456 0 -1 5410
box -4 -6 20 206
use FILL  SFILL44560x52100
timestamp 1596033377
transform -1 0 4472 0 -1 5410
box -4 -6 20 206
use FILL  SFILL44720x52100
timestamp 1596033377
transform -1 0 4488 0 -1 5410
box -4 -6 20 206
use AOI21X1  _4283_
timestamp 1596033377
transform -1 0 4696 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4417_
timestamp 1596033377
transform -1 0 4888 0 -1 5410
box -4 -6 196 206
use MUX2X1  _4205_
timestamp 1596033377
transform -1 0 4984 0 -1 5410
box -4 -6 100 206
use OAI21X1  _3770_
timestamp 1596033377
transform 1 0 4984 0 -1 5410
box -4 -6 68 206
use NAND2X1  _3769_
timestamp 1596033377
transform -1 0 5096 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4327_
timestamp 1596033377
transform -1 0 5288 0 -1 5410
box -4 -6 196 206
use OAI22X1  _4200_
timestamp 1596033377
transform 1 0 5288 0 -1 5410
box -4 -6 84 206
use OAI21X1  _4199_
timestamp 1596033377
transform -1 0 5432 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4322_
timestamp 1596033377
transform -1 0 5624 0 -1 5410
box -4 -6 196 206
use NAND2X1  _3759_
timestamp 1596033377
transform 1 0 5624 0 -1 5410
box -4 -6 52 206
use OAI21X1  _3760_
timestamp 1596033377
transform -1 0 5736 0 -1 5410
box -4 -6 68 206
use MUX2X1  _4197_
timestamp 1596033377
transform -1 0 5832 0 -1 5410
box -4 -6 100 206
use MUX2X1  _4019_
timestamp 1596033377
transform -1 0 5928 0 -1 5410
box -4 -6 100 206
use DFFPOSX1  _4386_
timestamp 1596033377
transform -1 0 6184 0 -1 5410
box -4 -6 196 206
use FILL  SFILL59280x52100
timestamp 1596033377
transform -1 0 5944 0 -1 5410
box -4 -6 20 206
use FILL  SFILL59440x52100
timestamp 1596033377
transform -1 0 5960 0 -1 5410
box -4 -6 20 206
use FILL  SFILL59600x52100
timestamp 1596033377
transform -1 0 5976 0 -1 5410
box -4 -6 20 206
use FILL  SFILL59760x52100
timestamp 1596033377
transform -1 0 5992 0 -1 5410
box -4 -6 20 206
use NOR2X1  _3826_
timestamp 1596033377
transform 1 0 6184 0 -1 5410
box -4 -6 52 206
use AOI21X1  _3827_
timestamp 1596033377
transform -1 0 6296 0 -1 5410
box -4 -6 68 206
use MUX2X1  _4252_
timestamp 1596033377
transform -1 0 6392 0 -1 5410
box -4 -6 100 206
use MUX2X1  _4074_
timestamp 1596033377
transform -1 0 6488 0 -1 5410
box -4 -6 100 206
use NAND2X1  _3793_
timestamp 1596033377
transform 1 0 6488 0 -1 5410
box -4 -6 52 206
use OAI21X1  _3794_
timestamp 1596033377
transform -1 0 6600 0 -1 5410
box -4 -6 68 206
use DFFPOSX1  _4354_
timestamp 1596033377
transform -1 0 6792 0 -1 5410
box -4 -6 196 206
use DFFPOSX1  _4391_
timestamp 1596033377
transform -1 0 6984 0 -1 5410
box -4 -6 196 206
use NOR2X1  _3836_
timestamp 1596033377
transform 1 0 6984 0 -1 5410
box -4 -6 52 206
use AOI21X1  _3837_
timestamp 1596033377
transform -1 0 7096 0 -1 5410
box -4 -6 68 206
use OAI21X1  _3804_
timestamp 1596033377
transform 1 0 7096 0 -1 5410
box -4 -6 68 206
use NAND2X1  _3803_
timestamp 1596033377
transform -1 0 7208 0 -1 5410
box -4 -6 52 206
use DFFPOSX1  _4359_
timestamp 1596033377
transform -1 0 7400 0 -1 5410
box -4 -6 196 206
<< labels >>
flabel metal4 s 2912 -10 2976 0 7 FreeSans 24 270 0 0 gnd
port 0 nsew
flabel metal4 s 1408 -10 1472 0 7 FreeSans 24 270 0 0 vdd
port 1 nsew
flabel metal2 s 3821 5457 3827 5463 3 FreeSans 24 90 0 0 adrs_bus[15]
port 2 nsew
flabel metal2 s 3501 5457 3507 5463 3 FreeSans 24 90 0 0 adrs_bus[14]
port 3 nsew
flabel metal2 s 3709 5457 3715 5463 3 FreeSans 24 90 0 0 adrs_bus[13]
port 4 nsew
flabel metal2 s 3677 5457 3683 5463 3 FreeSans 24 90 0 0 adrs_bus[12]
port 5 nsew
flabel metal2 s 2845 5457 2851 5463 3 FreeSans 24 90 0 0 adrs_bus[11]
port 6 nsew
flabel metal2 s 2797 5457 2803 5463 3 FreeSans 24 90 0 0 adrs_bus[10]
port 7 nsew
flabel metal2 s 3021 5457 3027 5463 3 FreeSans 24 90 0 0 adrs_bus[9]
port 8 nsew
flabel metal2 s 3469 5457 3475 5463 3 FreeSans 24 90 0 0 adrs_bus[8]
port 9 nsew
flabel metal2 s 3565 5457 3571 5463 3 FreeSans 24 90 0 0 adrs_bus[7]
port 10 nsew
flabel metal2 s 3165 -23 3171 -17 7 FreeSans 24 270 0 0 adrs_bus[6]
port 11 nsew
flabel metal2 s 3213 -23 3219 -17 7 FreeSans 24 270 0 0 adrs_bus[5]
port 12 nsew
flabel metal2 s 3437 5457 3443 5463 3 FreeSans 24 90 0 0 adrs_bus[4]
port 13 nsew
flabel metal2 s 3565 -23 3571 -17 7 FreeSans 24 270 0 0 adrs_bus[3]
port 14 nsew
flabel metal2 s 3117 -23 3123 -17 7 FreeSans 24 270 0 0 adrs_bus[2]
port 15 nsew
flabel metal2 s 3661 -23 3667 -17 7 FreeSans 24 270 0 0 adrs_bus[1]
port 16 nsew
flabel metal2 s 3501 -23 3507 -17 7 FreeSans 24 270 0 0 adrs_bus[0]
port 17 nsew
flabel metal3 s 7437 3317 7443 3323 3 FreeSans 24 0 0 0 clock
port 18 nsew
flabel metal2 s 4061 -23 4067 -17 7 FreeSans 24 270 0 0 data_in[15]
port 19 nsew
flabel metal2 s 3757 -23 3763 -17 7 FreeSans 24 270 0 0 data_in[14]
port 20 nsew
flabel metal2 s 4109 -23 4115 -17 7 FreeSans 24 270 0 0 data_in[13]
port 21 nsew
flabel metal2 s 4925 -23 4931 -17 7 FreeSans 24 270 0 0 data_in[12]
port 22 nsew
flabel metal2 s 5197 -23 5203 -17 7 FreeSans 24 270 0 0 data_in[11]
port 23 nsew
flabel metal2 s 5149 -23 5155 -17 7 FreeSans 24 270 0 0 data_in[10]
port 24 nsew
flabel metal2 s 5053 -23 5059 -17 7 FreeSans 24 270 0 0 data_in[9]
port 25 nsew
flabel metal2 s 4781 -23 4787 -17 7 FreeSans 24 270 0 0 data_in[8]
port 26 nsew
flabel metal2 s 4861 -23 4867 -17 7 FreeSans 24 270 0 0 data_in[7]
port 27 nsew
flabel metal2 s 4813 -23 4819 -17 7 FreeSans 24 270 0 0 data_in[6]
port 28 nsew
flabel metal2 s 4893 -23 4899 -17 7 FreeSans 24 270 0 0 data_in[5]
port 29 nsew
flabel metal2 s 4717 -23 4723 -17 7 FreeSans 24 270 0 0 data_in[4]
port 30 nsew
flabel metal2 s 4957 -23 4963 -17 7 FreeSans 24 270 0 0 data_in[3]
port 31 nsew
flabel metal2 s 5101 -23 5107 -17 7 FreeSans 24 270 0 0 data_in[2]
port 32 nsew
flabel metal2 s 3997 -23 4003 -17 7 FreeSans 24 270 0 0 data_in[1]
port 33 nsew
flabel metal2 s 4589 -23 4595 -17 7 FreeSans 24 270 0 0 data_in[0]
port 34 nsew
flabel metal2 s 3645 5457 3651 5463 3 FreeSans 24 90 0 0 data_out[15]
port 35 nsew
flabel metal3 s -35 4897 -29 4903 7 FreeSans 24 0 0 0 data_out[14]
port 36 nsew
flabel metal2 s 1245 5457 1251 5463 3 FreeSans 24 90 0 0 data_out[13]
port 37 nsew
flabel metal2 s 1533 5457 1539 5463 3 FreeSans 24 90 0 0 data_out[12]
port 38 nsew
flabel metal2 s 589 5457 595 5463 3 FreeSans 24 90 0 0 data_out[11]
port 39 nsew
flabel metal3 s -35 5297 -29 5303 7 FreeSans 24 0 0 0 data_out[10]
port 40 nsew
flabel metal2 s 2589 5457 2595 5463 3 FreeSans 24 90 0 0 data_out[9]
port 41 nsew
flabel metal2 s 2557 5457 2563 5463 3 FreeSans 24 90 0 0 data_out[8]
port 42 nsew
flabel metal2 s 2557 -23 2563 -17 7 FreeSans 24 270 0 0 data_out[7]
port 43 nsew
flabel metal2 s 3069 -23 3075 -17 7 FreeSans 24 270 0 0 data_out[6]
port 44 nsew
flabel metal2 s 2509 -23 2515 -17 7 FreeSans 24 270 0 0 data_out[5]
port 45 nsew
flabel metal2 s 2221 -23 2227 -17 7 FreeSans 24 270 0 0 data_out[4]
port 46 nsew
flabel metal3 s -35 1097 -29 1103 7 FreeSans 24 0 0 0 data_out[3]
port 47 nsew
flabel metal3 s -35 897 -29 903 7 FreeSans 24 0 0 0 data_out[2]
port 48 nsew
flabel metal2 s 717 -23 723 -17 7 FreeSans 24 270 0 0 data_out[1]
port 49 nsew
flabel metal2 s 541 -23 547 -17 7 FreeSans 24 270 0 0 data_out[0]
port 50 nsew
flabel metal2 s 3693 -23 3699 -17 7 FreeSans 24 270 0 0 mem_rd
port 51 nsew
flabel metal2 s 4509 -23 4515 -17 7 FreeSans 24 270 0 0 mem_wr
port 52 nsew
flabel metal2 s 3613 5457 3619 5463 3 FreeSans 24 90 0 0 reset
port 53 nsew
<< end >>
